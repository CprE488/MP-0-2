XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3�m�C�hǂ�"rϱS�ō.nC��8&� 0l7����er���ϳ��Ҧ|���y��P�,<����;�qI]�(
;���c|-.xOљw�`m#N{Q���n�cTU%��OCyeK�-k����N�l�Db�:a�jw��J��,%{a�DZ��^����\���f���^@um�zDB�B�{_�f5�ˠ��(���g-�

����B�V����}��<N��A0ʮc�6KKJ$J(u���/�֌�0�Ɣ ���J��~�)v�Y� �cm�ԑ�w�ǊǚA),B�&nH�X���dd( �Gཱྀ����)&�����`\[�q����x�(���?>d��R�(��0l��dǕ���5��iOuvw�mY*�宊���c?�'��Y;ܣ�]����B�i�Kps�9��z0���#b�({�0��fT>��^Kr�v��ɔ������ONhc������n"!��Ͷ�3������Ը��J=Tw7Pߦ&�D]��o~��X��T������*t���:d��s}��mv�L�����=*�[In\��������%v�5j1�8��r]��q�r�ZN@ݒY��Ul�6^��*� ��t܁��P�k�k��t��8�{�y��~I��PbO+C�8��H���:{�4����5��h��1K��s.���C#u3�1�z�Y�5��y�-%�l��A��~}��3:�.��~\0���)�'��B�JdQ��N&��%_Ō��(�2F]���$�؝SY8XlxVHYEB    fa00    2040)d�;
��<
K�ހ����� ��W��u��<�SJ��S])�
��BG'ݿX\\-R��iϛv$Sf7�7:���
�򸒓�;��z�����L!�6&���C��T��'��?������w�(P#�Ib�&��ߋ@-�����}����}l�}�]�;B_C�l��)p޷Ef-���˿�Y��G%;�h��͂����O�
��?+��OX��q���g����]��i�tm2�wc�3 ��v��K|��MJ����z������)�jU�WME���W�7Ji�f�ų�b��@,��S{@Ǜh��k��eoix�k'U���_�M�0��'��ˮ��[�����J�_l�Ab��V܎�C��Rq��bWv������q�ʲ[ݙ��l�Γ�^9]����v��|�>�AX�����|Ι�)�k��eI�鷎�&�>��5�����"F�pl���fe|�e9�O�|���p�P9����W@��\�[���'X4S���D��w�G��,S��w���cǷ1OM[��r���B2���F�~��D[�Zk�[�Z*�hW�#�����1z�l�<D�����Bx��ʴe8�ϭ�x ����i���BU�n�%;;�l���l-�� A�Ŧ�&���ro�������7��-��wb�m~���h���&7��e��B4�!r�}J��%I��QT=UU7���A�h�W��zH�u�O�C&+������W?Bo�1jVB m�P$�uJsQ[v� ?�A�����䢗q�a��Nx�u�����G���z��)���"��d/!�(�nfPW<�T�)��[�x2Ӳ�"� �x<Va��J�G�d ���`���]�[��(���F���:;�nfa5
��hH���Ӝ7�So�
Al�2�(�He�ns+�O5ϟ�����A�Invȑ'�?Sy$�@��vpǓ���*u2� s�6�C��h��O�"�b`l��vt��<H��m����5B<ۃ��E�M7H+FO{С(��!��iR|0�úET��O`*�#x�-{�Ҟ�p�(ż ���zxf��:7,����(L�%�?�B��_%"^նW����b��&h�
����Tؼ���)��P��9{�d¹�R�XZ��TL�>�u��)ƣ+5]z�?�۱h�G^tݱ�ކI�z|�����x�M�T�5�f�F,���G��#��~1�Lj�����4 Ek*d��%�[ۣFC2h'G-��~o��˦JC_�a/O�e:��I-���Z�QUP�Ux�X���|��1����\�g���IsPX~}�]�v�U	��>gɶ�66d� �<hKw��l���?s�7.�i&)n,@⑍v"&��Eq:��l�ߥ���CTqd"���á��]�cn�fhN�0�/�:����H�wa����x�@��xjd�,����"��%��k=�����5^7$�B7�F�zWm2En�!v�k���5�������kS���Ӧ*�l����݇��-��Lz��B?Ě�>��$B�h�PH6i
�b@4�*䑌����	�R�`�в-|dGk�I$+i�y;��Gs2S�o�z�7��R��?���Y���RZ��V�����?U���M��xX�t�5���q����p�c�َ�m~[r�T����{����H2�ڽ6��{�v�_��ΰR��4Y������ˠ���'�pR��i\E�����!E��g����Rub�w'�6��3��� }�҂�@]2�7L`Zϖ��
���H���0�ҝE~5���%�{joܶw����m����r+	�<�ӾDt��dUb��[v���f�a)^���3�U���p��D�{�4M<��)��)��'[
v��m�%�қLrGl��WL?Q��RUI`)J#>Mq	�I0�Y�k����A�u�E���wz�	���e�ެ��'
��]��Xҍ�+�����ҩ:P�8'�Smv�b�V�����g�=N��8]���OJ�xQ"Ɖ�5��:���!���(u�^4+9�&���ZaE�QDƭ���������Hbٙ�XL~4��O��������靈n&��~�1`�K�ɪ��1V�y��VXV��o���),�i�ss-��w��;�4j��FV���˦)f�<D-����|ס�-��}��4^��2]��
�m}��R~�U~ôe��A^}�cN�dJ �
Ŧ�@�T�s�屛��gu; ��<R!���A������e�⩻ٓ�ֶ�����]�}G[�w�hA�G�&�Z�*mc&3'�h��b�,��x�Pz�8*�����=�TWj��T���N�ub�B/ֳ���*|���P���M��OR�9P��uTMQ�%�3}X(��u��a�]���=Q���׏�B���"`��c璝��:s	̟b_W�b�o�_c�rl�S�S�4l�lKR�uĵ���<7�l��t1���^h��n,R��m�ąV����!C�����:+�e�b0����N�-��)g��	�����z�ʞ�߰%W&�#��U=x���\D�R�+��?T�l^��v捬�=���[�b��2������6���L�h>==;��Tq��&���QH�e���A�AX)�U�>O9e�����i��o�@S��U�K���["@aO�~{I]���1GʯT���8��Ĥ@�BB����d����4���:39�� �1��_��
���no�p�!���o؃��j'3�n�Ը_3�̐ֵNl��a��Z�ug���d�Ţ�T���&�̈́��Oo�K�VAs�5fG�3��k��}[�pL��{� c��T�GH�9��I<(���_ҊXu�5Q�#��X��*���9<��R��^�Wdբ	��/��D��:�cFF��3����n��~Yߗ@B1 �pM�R ϳ�	%��n��
�W A���9����ɺJ�����pM�:��E*�\lyx�1�6.8�h�A��i����_k��x�w�"�9���&1�0$���]�����^�E�\�\a�卛��*^�f�&3�gy6D� BJ��p���I5G�<�J8Y_^��58}Q�Q�,:��^�!Y�d���ݝ�fHUR��G��N{#��믌��i�G�{Ȯ�
Rҙ�%�V���oQRQs,����f-��$*�S����9��M/�_竟��j���� T8��m7O�
�)�ʫ!���:���m8�5$rVݖe?��v�L�U�y�r,�T��#�%�iq���6�����G��"A30=~��"21��&$��+��h��xU�f�%�}����Ȁ��Dz�'挄ȟ��w?@1����aE��[�Ur����T֐����j����I�w=!�[��^sДkT��5�x��ޖ l�?i�H�MȺKeX�С܉ ��'�$�ܬ0V=sLFϔA˰h����M�(y��-�]��g���5wȱ��g`�+�_t��%I�vmH�Ć#ܘ��s���o��z5T�{`HJ.J��+�IQ�~)ތ�0��Es����r�Ќ�F7=��|�R�vB���^\�|���v@#�hS���:�h p?��.4_%�N?�a�\@5 t���d	ɴɰe�u*�5��6��M��nt��/HU���^V9[�����xgqf4C��ŐT�1t�=�6�������gW�9�UJxЫ���!2���8�B���%ϚB��'�b[�[�RNW)|{��j{"T��쐝��/���k���1N7S^��ǅ(�]�?�P�j���y��C4���6�#ր ��L��|lp�J�3'�`L*Q-hE6I�Q��HmR5�H����X��1!�j�5B�	^ u!��7�(%�f7E!@��p̎�U�܎ia<��&wšA�� ��K�x9����߷A}^�󶩲	�]�\�Ӟ�Kn�����X�1{q��J��t�)�����(�+��P�b�붴ɼW��F;TT�+�A��3p�	"ڞ��2�Lc"�������-��M��y�Yj�mc���tIO�D�ch�x��1�x(;�Ř5M��I�MU}��%�>.�O�+;u�D������%u�����}1V���O��=�,2H����/+�R�����I;k��T�މ�2�r5�X�;=N*M���w��{R�Q�����0n;rO��:Hes���%3}ۻ� �����TƘ��R.u��4��a)_�Ct��WU�m���%�x��O�F�c]K ���t�ڋ�-�P�wMM�35�rDZ���>��ia�Ǹ��`c��t��kɪ�K�0̋Ķ �3]V�
���>�V[��ӿ�G$��Қ���V�{��������5Mdb����45�![?�aj��,t�.	*;����e:�Ɋ���9�AFH�����7F\q(0Y!�2�7�D�.�0n�웽r}���==�O�bY�Z%�)D�|�v�ϰ����w��
o���p��t���J`o�f�ޅ?�Hx�eK.��걕B��+YvK���tG��ń�q��a=n4�fc�uX��IRw�w�pr$�M���Vp*/���bs�|7딤���B���M������ϞV��g�l��B�����>(�ӼԤ�����n�����.^ܦ\ݎ���7%�&$#���?��^�e��o\�f��('��Z��D���o�s1d�E㭋���mf���-��~n"q���0#�&��l|5��f ���(�"-ʖ�����@�u����RM�����`D��H0O6���z�ߋ0�/F	���ϳ�_	ؠ��쎕 AO�Y�D%y ���&���~_�َ6�:}]O_�UYY�Ko9��:��~'���ˠ���8!_pb Y?������O[yf�|{NB�*�G�s�ˑ����g��_(����#�������:����ƅ�
M�_/�2yů�?��*
�Ұ����\�Fn�f�-d��Ҹ���)���v����r��g���X��z����i;�sn�A��yb�TC�8������DN��f�Z�G��Z ��!L�Ig�֗���Y,k��J��q}i�j�PMŻr�D\E��~^F�0i;,l$2ēO}!�'n�9�B����C����O�F�x�����:���Hx�K$�BǷ���m-K1�I���_u�egd�����)t�y�aA؇̿h��Gb[i*K}��B�������B?sm%���vv!�Bh��>rn�0#���m9,9��y�ePn�2���(:�{�zF�'kEy����R������;�p�a�zr#�!)e_u�A��q*Ļ�z�$w5�?���_� ��r�C�����1���_@�d����zۡyfD�<�j�jF�p���"b1 [��-��?Ǟ��AGc�qW������[7�;��`���@�h�����d�I�F����_/[L�W-��ŀ��8T��q����ܘ�=t��y�l���=�+oI��hᮺ��ֲ3�Qi� ��`#�џRѣ�MKTYWJ[]�G`��Rᐊ���w?�y<��y����v����Ō�4Q �O���q��m`|j���{L�#�ݠ��mu�fX������LGqOh&�l>���n5���tlPH���S�Q�D=<���٦���lٔ@y��O�c��@J	Z�Q��$I*��&���_�x��_� �k�|�	J
B�-��Bֻ��L��X_N�o�;i\"��ů\=m������~J�p+�����fPy�Ć�TA�K��k��,��zT����(��FG�q`iN���QU���X3c��羧m8��* ,���ݞ���3p���_�T��E��[�lR\�z�.җ��8d������v��9�����w`������Y\�u���>GMYc��:��p�e�I9�7e��g�QL��۸�"��t�'� ��7y-�6��T�r#��wß<� ���?�z��_�[VI�FM����^����j4�Dj��wA=�l+Ng�L�S���rN����݀�y��&�G�3A	;@��_��$�� �Իq����ąy��4�t&]������|�����U�O�x�m2��g��~�Q���/��z�(N�Ya+����p�ۖ\ú�J�8_��|���4�;�l���2��=S�G�R�vfq�ЪM����)����cQ�*qj��9�]�ǙQ4eE�ӽ-�7F�L�/��M�[2��J\e�
�8���j^�W��Q��$|����½�#|]��Ah�e�O�C?�`T�O>KB��-:���3�:����l�%7����g�1�Um�����r���O���m�!��·!8}��S�H�@0��W��>������!�OɃ�6o�7�;���3��%��~�ͭu2���Z��c��%��	r0����p��EC�[/*�ڧ����i�?wyz���*_Z���To�����4���C����ڑ��j��{=h�:��h�^v9�Ԭ�y�׿P�G���,�~u(���h��}�ί"�I�dn���;�J{s#,:�FsóIa/[��߆�oT�R_�U��m�����2C8ѳ�{���x�s:�1P1|Ѹ��=����.P6��'��L? E{M}x�M[��+B������^�~������&���$�w�w�p���?
�hׄ7T�K�
ы=��0�q�(���������r�Uo��-����<5<�;��6�' ��5�L՟�w�RY��G��K�P��qs]�9�ft�]	�-q�������DT-�m+���m��Q�ڸS������0v�]Ye(yh����[��H��%
�[�(�!C#�Ȁk��t���	�����ֹ���F���D��|�l��tR� M\�Dv��s,�ԎLfX��cT�[2�|g���4�R��q�1:�6]¦�F�O�W}������w,�䇞c�����Ʒ����K]	���G����|4n�l5���h�r�KG��k�J�b�7�U��V��0ŞOA�Q�!���P؎a��]�y��K�O��$*��@o+�*s�>h�d�Kb��7���x�7�Iư�Q%�h�d�u�[�C���*T=ޛ������FT$�k�v��#��,�s��N.�Aߎ�������C�m�|6�x9�].�4UL&����-Y��(���9����H"��+9|9Y%��p�eձ������4��D�/�q@v,��JQy�X����gA���v&V%|Y�q����d�E�����(�%�84|�Rx��gZ�D�4���=	� �[�}$�q��{Pb�^�Yz������rOI�qm��;0ųM��6�-�Ǫ�k�!Ӓo�J��9�T%��}о�)�ŹF��.[c�	��OܓL�ӧc����܀�f�� i8S� ̶����KbV\�Qv�:�E�t�����y��������ɼ��7�?�+���9Ƈ�..���	��$��Wߓ�=ڮ�n� �Ztvo_���K�C 9/���������(�m�ѺR�w��;�J1YnHM0|��S [��˷�PC(�~�=�7��^&_%L�e����<����Uv� Ӿ�Il�
�+�S�[�>��{��5J�cI�H\�������w�7�UGn��r�tK���
��/��Y���&�i��% �b�5H˷�=4z�Fe�W��k>�;;��q�u�n���F�]��(M�4�*K@�/��e�͚#�|��Q�������B�3ٲ8���U|{k�W�nM��ʪ�� +�a����}%�%� ���,O�����K��n(�Z�ִiDD!��������A���UE��LD	�^�x�fx;Z;�&]:7iއ�wo
j|K0����/M#dm�����:v�l6�,?�r��d|��:Rv4#�W�7���[�x,^����'�ie���_㔘�Z����#�?�o��/�
���"�m��У�zGبyH3��3�\��pDR��l���"����h��X{��3���<�R��	
��(�Z�w�|�'"�r�ͅ�,���z?[�Ic{�a�(�pX�AIZ�)u(׍F.�
�����}�CU�b�v�38���Z�^~K�l,���ر�[+E�������B�m̀<�_���[�f2;]�K�3��e�Ɩd`�XlxVHYEB    4f62     b50n U�����d٨P�xu�S�K�#�z���n�e%��<w�.TXDlW[��2�5_-${	S׬�Ρ�^�`�p�fONqxJ��D~��ќ�4�z�<�;w��w^���S� <�)�e�ܾ}>�_�!g�S4��O��w�I��3=.lꑘ�eG�C��e)H��h�9qc��N��4�X�7eie��شif�����ssZDd�7􏥝V�Ii1�xZ�V�	�Z8R[@�"&�q:@q��׳.h`a�xu��_4�4K��o���l\��x�:2�v5V5*�J�"���,�1
��3j��k����"�ۋ�5��|W߶Aoh��x����~��
�pV��N�λ?�J٬��H|Gއ�e G�����i?ы�i�L�7�c"��6Ʃ��= Y&	�m$"m�
~
�^����k��&��_4��Y�\ե�2&��O"#*Ul$7�9�Ӯ8Ic?��cy���/L:=ǫ�����KK�b85^�����#�@�G�{"�ؘ_xG�3��u1ɩ��ӛxa0?�ʏ�3��~�M���sj\�Fү=�� O D���9�("9�_�F(7���nυŃ�D7��n����c�z	�Fb� �6\wΤJ��keߞ��v!�1�!&O�VPb�>d����EV�n�ؕ��/�\��[��8�\������G�&��Z9�A�`�+�S~!-�����)\�]H�L?^xp�/� =��b��^	��"p<��
`n��G�]�ٍ�Tv1��i�m��/�l��&���b%��+�0�gEoU���>S9�z�.ċ*�!F��	�W�>���bc�������Q�&e�hW�Ճ̓I"��$n*$V�&#}{�k~aAK�w{���"|��)�`����"e�����f��� �� ��v��SԔt"����d��*s�%^�%f(T��sb�&'�����������N̈́�`���r�}��A��vL��OfJ��e�Ge����@"'�A| Z�6!(��Rv���8P�P�l�d��$ȝ��v�T<R���˝T�J��E�g^�#z����H{��K�Op,6ds��i�0]@���(��	;j�;��L�j��ה�=�$Ry���+PAj�y�SL	�"��F�Lp���;dӃa	�Lk��N��C�ɪ�L�5�x7A��S��j�z4l#I�`S�9(,�ut)�wg�z�d'�s�/[\K|@�_Ÿ�U�P�i6���OdRd�*(��:G5��+�|�w��|���:E�AP�B'�k��ؾDj�OQ��'R��SaB�NC�5Vfګ[��+��+ܧ��\B�UEG���˂K�x�"���p[z����ұ|�5�ص�>��y�hh/�q�Hd�;8�����X�ɡ��������x��%w)������R�>5[�+-j@	��"�&P��E��Kԏ�G2F�-�(0)�M>��>W6��y��_��3Pf��p���G���´��.�§H��<��� ������`O0�*�Ē�#�Fh����g�Μ���e/z:���Z���f�=^2Ӝ�Ke4��&�� ~��Kqp΋ċj�u�}�@t��H�=f��}��#!�S�����%����0)�wwP^\T3��F�/ X�-�������1̸N��U�̑���xeA}�(/A�*JK�W~��yq����i{� �$�C�0��o��0�Qyq��ܚ��Ga��(�V���a42N#i��~�v�3�w������(�C������:��{8L��.͹���D� �q�+��C#��ه�*x� �<�#|"}|���?�܁)S�ЍCa�t���r�'�W6>W�i��u��#��f���sn-��=�����K���p�9��͑��^o�^&�� �Z?pV��!<��[ѷ���_�ޗ�A�w6������3_�����9� �K���!r��a�
Y?z	_gC�?I��3�V�|�L.	<�틡���CksΙl�6�������W�g6lj%���� ��p���$|��3\Q}mj�y��Ƿ�@A������Y�wV३�=�M�ꏞ �����,�8���k�֗������`�)��Xx-���Ʉ{��Ϩq�3�ԯ-��ޤ�9��=�$q�7ϲg~�g��YA`̇w��Ps&k6�Y�?� ������x���2l5h!1�����,��ue�m��q��O�b�$��s�S��\�"�����pQ�j9�1�gEapI[�!���.�����!���Y�`��i�L��}L���Ư�5<�$ o�� ��.�(s��&�*K��ړ�O9
�q��F�g�q#���n��ľ����ovt�p�:� ?��5�_������r��5��?��\;�:����o���ݎd�]��߽v���k�E�`::�/����$�Dc�3ia�7��D1�����6��4f��u ��rx5u8����%&��)d�j\�n�]f���^r��.�'�����JRM �ͮ��ҟ�W��$he�IM�tp���R��Osh��4qf?�T�oF{��y{Իs�sh�\yw*p	b�~_[`i�X��A�e��IV�P��V���~��$�+PXu֚��DCon���?����TᗶQ�pi�2��նN�!�,Ps�I��D�]�4����;��cT����(���z�?{��y�<�����"3�5G��[�I�G�)���W�D��_��Q$�!ܭ;�#����O�&21�q�B��0@x���t����Ә���h��y�:�B�@�c�����p#@Y�6�OTu~��qy����k�FǇ�=@��:O
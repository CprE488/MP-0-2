XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����#�ܭ��S������dd������}٠JZ!H�غ�r�)��3��WwA~����������.��c��H}�L�}ɤ>g��
�Q��A�+:�!4k�Z����np�1��Ju����'O�|�<�b�زr�˕�rm�\� D�6�m�5�)́1T2g��ԦJ5��c�5WD�6�҈��2�K�)�\��7GkIuBP���w����	<ٝ�%�J�p��ai�l�(Q���v2�$�Y�u��**�$�h=�#%Ӵ�������d��t��v;�^|���|�,�;k����ԭ���a��u*��͗����&ꌩ�~N�A��E�!�m�B�$I�:S�>��!�HM�ǥG}IO��Ţa�Q�]����I��L���Ϝ����.IƖ�=�-��K��͕�0��U��z���/��8{���R`�zZ��N��ѹ71��tJg������VL*Q�>"�R|v� 8?ê�(�~D����~�����g�V�ֲw�j�}�O]����.ءG.9�ɿa��Y�I�[]��u�/.������9�,c ��q[�s|��΍�(bfĖa
�d� ��5,f%Q5W��OeB��I�c�����Y��5I��\�G�����ϛ�����y�`���	���m;Xʼ5��Yf�	Id�<,-4�#���({�����j�ץ�ݹ1�� �0�1���уb])��c��\+��x�#�B����(Ѩ}�Ϡ���GK���w[w�ST��XlxVHYEB    3fdc    1160�T��Ā�J���P�S���80���ҷ\�H���VW>Ӫ��."�0��j��ϧ[���Ys:RZ&e=�l���碀$�"=���m~6p��h�CT�E�/D��-��f5�|U��t�啩�п�"ޑnQLL�4 N��wV�Js`�K��ߩB$�������u�U5��'����Y���o�l�8~r��Q�e"��h87��z���F^���*4�D�����s^0�ߋ)Ѝ�7�S.'����6f��E��j5d?Nj�<E�ۚj@�k\�y��|ҊM .k��4��z*�Ȑt��S�ְ]ON4�@���~��o��<��ĸѰn�\t�ҘhU��5 ��N�sv�b{���v�ZWݝ����\g�@������F�ت�6�}�{ޗ&�XT�*U����V���ᔡ=��)����/�f�"��ՠ���2@+��˟�T4��	&p�hsoO�0���f�9*�e��U� 9$z���R,����I�`�Z?���"	O|�(������"e,�����X+�mq�G��ISBǾ�m�`b�	������e	�dr�t?3m5q_�����IMHD<]iٰI���� ~�`-L�ˡn����?w�p
'xl�8h�;��a�7�Ct5��lM`���u�Z��3�U��s��)��R����(<����w�>��%�ě?�Ţ�|żY�x>t�|�3D����q$�\ɧy�Fe�s��n�s�=�柱��d�U�+Ј:>;cO��V����܆���;d�ܑy��>-o�"<��8���m�I:�ۑ�M�[��LpŴ�/���(����U}��:����%�tO~2V$�Lh����5������/u��������6(�o]آqR�����q/Ċ�˧�%5�n�,$�=*�Z�`Ʋ~�io8#(��+SZ�oMRc��W��b�6v׽w ���RR�t- ��,���9}XD{�̲� Lb����Cܛ�t])��+�'� ��] iQHV>%�HmJ���W�!F�Y	��	BW����˂c�S��O�ؤ����; j�Y柺(J� S/�X��Av�����^��$�jQ2���cT�0�zre^�J߼�K_��҅��y�����*.A�~X�@K���x��K��?%l��|��f3̾G�*:n�k��e��?Kj���Q�V�kɒ0p�0M�`GX2`w�h%��ݩ
��u������W��K��J {NSY2�s/�v���G94swpv�9��C�fɂ�2�Y�l�iӪ"�?�^�Guׅh#�2�	��J���&�O�]��y$܎������h����2����`0�K7/��-}�s�*��g��y�9`Jq��}f��ȬŵW���\�5μ�^�7��XS�ЫoL�ֳk�i4��X1�w�^-�f�Hr��M=���I�$��	���H!�En���9�^�ƅ,�=�O�<�K�dҜz���T�o0���I�PX��C>(��5O笒*dM���eE"�܉���k���&��6���ۜ^�V�$�_�\.Qý�+�a����
}W?��s���2�.-��k.�G�lG3:2�; ���"/��%���뮂��QP��i@�E�uw����l���<0�i���A�N1��߱��Q��A��[]���G��Z-l�Xt�Љ2�^�U�T���a��"���ί�]U��M�!+�)�k0����C~ݽ����/w�L����AR��0��M�#»�&.G�v��3#Qhٌ��F4��h���_.�Q�1�j��d�DFR������;I^�x���4���y�O�c-�f�5t� =%�F�p�+���2����:I��d�7�abI���큰,���7��R�[Vg/\�м@�h��b�����ݧ�G�	���Ι�Vw��@���-DDs�DT����^lC��e�jj���pb�Y8W�1�PZ�[�>97 �>F0���Ù���u�����0�I�莟{�ܡ�V�Cf�Czp>����@^P��$���:��xA��m~�n 7�s�>a3^��.��z�7�4Ms���ƺ~�J��}��ys (�jk����7�)8�l�DS�𢯟�h����(ޥ�N�\�O@M|��9	xF�=H:�,�4�UEF����A�ک�y[ �,Hn��r~`�>(<�
��{{2�����M�
N�֫O�X')��T��am����&LT�$C!Z���-�t���cl�R�D"p���+3|���^u���=��͂oC$"�FiM'������x�-5>���r��OD���<6��D D�5M�%��Î!���	�;�p)S�7 h��x��v�87������K����g}�bF�u,c�TJ�\-ϟ��I������["�l�;���qUɣo�7�:���ޥ�+[������@����9mZ�<��;��|���'�!-s��;c�jQU�vF��Ԍ��Y~����M,m��f�-�p]�ʆ���������Z#a�\_�Բ�#
h����u�H�T�3XR��#�Wٗ�A�KR9�&Μ���B�=zD�l�N7}3���bIP|�󝒃�8��2/A̫�Amk�a���q�o��cD&�P���,��~C�z�ˡ@�}��1 *�-���YF�F��r΀"�%i)J���EЃ��>R�4����f��n8&W���=����؁G��C̜-���ԩRr�h�j�	-ƨf���)1�wr�mw��Sy5
3�����%�I��q��;���m/� ����ߪ�@4���*�0ϡ��q��@6-?�	]��'��{��[�;-g�z�	�Dz�}�0�a�-��AE�7
Ʌt��>n򊡵�73����l��\)��`��p���W���k�	#(���6��W��n��g�՜��amٹ*��l�A}z�� ����ݕ��e����P���pC�p��T{��E�������{��d�%Ae�HS�����[t�I<Re�l�և�݁�8=�3��{�4�d,Z�j؈y���ՠR	Yds�=�Ck��ۃ�j
X��q�����2�҄y�xs��g�h�6����3(��Sd��0#��K�O��V��R��^�u@%V���i����*� pe\�,��|�{�]U�ta���H��ϸ5�`�����"� {�-�u�7��+�E/��Z�P��gG[�5�/��b07�bV����[t�7Nf�&@]��� ��h��N��j�,C���3��5�m�X�����A���W�Տ��l!x��"4
�a������԰�~J��#}^�t���Hf�m@��<����a�u�6���r�A/�bp08%g�����%��`��9p;��2j�[V:=�2J�]מ�y��I��,a,T��ŴcX?�1a@�wfx'�#�j�Ji;�M+g6����|�t0H��%=�mO�}�ۯ�e>�Q���v�!Q���~ߓ*��Ȑeݭut�� ��j Z>�fk�n�� Ik�
�����	�3�Q�Q�������U�����靳�Ր��k�Ц�#va�Gy!��YgV�rC�[5�{}dۦz�x���<l�]��=�����f�~JO������1 yJ�(��%�Zi�"z��]�E����6,!��X
���O�X3O)RV��փ�*�.rY4�!�mz^+q2�T�(s�l9�IC�Pd���h?�^�����$�=����F�@�M�4gJ���N�j���$jJ)6�L9�g�2EJIu�O�Q'�y:#��8�)���9"�ឤ�:�N��҄/�<.�Fo\�w�o����1 ��7`���iJ0��:������'f�LC���t���]�sW�c�G	.nD��c'z&!'P�� ���7Ǌnb�CW�84N�����ձ�n�?� x�"�ל{����#���|�cT����w#�c��"?�i�^�{s+d;r�{ ���H<�~5Du��5�}x�.��Ku�SC��EB��M-cR�C;s�,S��D;�����??3���	 �p�D"����,����g���(����� I�����*"ލ8!�/ͨiusڶ-4�����'�!o xR�ocP�;���æ�Zz)ٔ��a{��L�M�J7�����?@4{�F�rWr9�B����c453qX��S�/�g`�9�����%�a�Hޙ�UD:cc�b3��O��4$�Q�)gR2���J_&���w��ON
�Mb��hU�Y�|�J�-�}.L�	-�N	x��Y'97�������ט���ba�ERI�$��z��f"�O�2n�0���֤4�^Q�3L���K�=��M��˻Z8��Iw���(�o��O�IM.�����WAO�82X,#j�ʹs\krL�.�R�D���&�Q���>H��Q�"GG���/�bx�o3G6�w�+�	�
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+HO���Y�o�����PE����n������]���w.p�B�1��A��ǡy�\���I���WȾ��:�.�,��ߧ�|�m���58����z���w�Yg�̡f�@���5��c���olް�UY\ĄG��j�ⲇ���"K��8�Q��8���W�=�׮�U	z��~<����5��Z��ܶP��D��iI|�xZ���n�;C���$�*��,��P=P���[�Rs�L
~�o ��Fb�Wh.	���A��#�K�1o䝵c��UXlQ�ǿ��q�0@:����r=�@&����<!f��j���"�-��T�֣p��8��>Dƛ^�eCi��ə^V����gC�9 a��0�Wv��{����˟`��fT�J+ci/� ��g���V^�`�w��,\�@.`�w�v�p�-�3(�MXU`,�(���2
�^G;�*�N�̘�"�TSlP��I'R��c�D���j�ҕ�[0؁���Z�$:N��T�tb}�Zj���� X
�������[�Ŕ��tR�#tS���k"��{��O�Vw�y�|�I�p�h>�/���px��<`��th�0��8���Z��ƴT6@�<�>w��:�C��V��5�c��Ra�Ï�u��G��kQ����R�`�0_/���첑p��;a�.BdJ~?��&M��q�`���p8��癏Vb��Y�y�Y�d�,��M��s��k�9�Б?��Q8Y��Bv�zi���XlxVHYEB    dd8f    2160�T ��r�G�^!JA�z�u�:`� (�Wkbh�?�2����s��q�A��C6�U �'��S�2�G��1�!�#� ��P�_CZ%�����F|7�`x2<EXn� ��2(nD���|M��6��}���ꪯ������5
S�RB�^��������Y5}����ExKMo����}�Jb�On��M/l�0�ʵC|����X��ʒ�>\�_��m�YP�u)��%�ˆ�͠8Z
㏢�ǝ�n���hN8Q%?�a��H;gn��0�~G�=���?s
ݘ��ton�+
�)�EϢ������g����D\<�JY�q_P�*���1ONVD`���W�JG���GΣN��@j�n�%�)(�K�.�	c�s�$� ����R <t̏�nLl��	͜Ҹ��:gL?A���o��W�{�lBG��
�ڃ��_k;��LE�=����u�9N��{���V9���4~h�u2�	��;������#�;[�`�=+�`,|�Z���tBޘ��U�\���>��-^�ގ:+P���U�-����J���f��AȤU�]�dF`��
���-@y U3$�C��$��@%]b��U�M��K.Dtn����� :� �n�y�1����z�_-��d"���!@S�t������o<�D�W�[u�̢�ZmU@[K��q/}��&�D,���\���� ��]^�H�[�� ���S�)[}����Cu ;B��?^?�Ͷ��g���*�Ȧ�F�r{��0e�&s���Os��2x�@���[N�����*=��"u��.	�w���D"^�
ݱWlޝ�b��9�ꆽ-�S�+|�Ｃ�y��7�;8}�R{�`�l&�p'��x����v���a^�_�k1�j��+�B��
Ƈ������|�(c�8��C:��Fյ�ٓ@�
�����Iބ;��;��<�;J�Q3���$��e�H�`�^5F/��ʖ�qk�'&�	t*H&��?���s zS� UL�y׉.��Q��3z7;��o����s��dH�� �^�Y�p	��cE��2��N#\������`��g��&#��~�!+b<��ł�������C�=��sn�Z���ک/�P�v�Zx�W����âc�z@$J
�)e����A3okm�H�q;�>��W�KlXƚ�'�ă�U(�5,�9||�(	�U*��r�~\l���=�!�/z��"�`�B�du� oOjg��B��3}�(�aoQ|c~�/�!-V�\������Bڷ�Cvj���1�^�H�C�"��*`��,4�,kE?���&d�;_��1���kyu��xa��~�mf�n4��䗖Tʿ���$��0ҵ�~��-��$�1���X�O��vN���Cx��k+�j�t�S�"�)��]��dq�PN�ro�3c�ݻ���,
O�	I|ؽ6pk3�0Eݢ,��P���sу��ݤ� 2̤�-Q�6��2TF��\�a�v�������h�aj�$n4-#��Y-*B5t��8���S�����ˈ��-4r�;�����d(��| �� �P��A��b�4Ζ�0Tg*��p.������\PH|��ꪯU+�q�tx�ؘ�mH՚��ؽ��3qhBԄ�b\>���ȱ��ys�qd����$V����V*�èʁ��H���3���G1⸦ǀ`��L��Ys���9i#.|�v���gh��@z=0kg�}VƊ`�8�m���4��`q�|%�ku���6�ކ�%�9]y�Y��l�w^�;�������������
��`���V
�G�܍q��Ξ����q]K%��"���f$J�B�a԰S��Tn���%7��ƾ��Pp����bBi��F�)��2{d��G$�����J�����;{�eSn ��\R񕂫��E��4b��m{Ws�i�2��{��1���@�v#�v��䤞���#�h½��E�Ga��rz����ҳ�����0J�q+��u��/�1B�P��FE��J��.��l�����+ٟ��p��)��T���z\Y��J��U
�t@�4ET�"X��q}>�-e�A9��2��ǎ���>cNTk�����1	1&��J�ȼf�{j�� ��2l�Za�m�Cu�a3T�wyzq�ȣ+XX�e�����p	Р���F^�PB^�N���'t��EDw�V������N����Av��G�
V=�p���$2�^5�,)����"�S�+հ9.��b�klS��Rvl������M�W���z3,��9<NEөj'xJv�*��)�x���m*^��I��m>�~Q����ЭP�!���
�w@|5�B0U�����A�%yԩm��qU�2���`k�����.=Gj.��$���s���[4�ѯF���t��ry5��7��c�" �T/�WX��j�	b�e�X�o��S��p3hv��xn�ۂG��sS�,�SӭI���X����
�����Q#V����2j��v�!��{6�H2�¢fE/'d2F�'쫻�K)a`4�
��`���~����r��Ȓ1���.�8�RA��#+!	u�U\�٣L�H��zkc��Ze13fN���XH��2!�,����kD�P| �<=L��D�
rl:�$y��AY�������i�ҋ�4ɢ�&Qx?��$�왍�h:�sQm��~O�^Gl3E���!��YG q8�����v������(�C]�=l�#f�q*��n�:��,jْa/c����C�7�����O���;�FQc=b��[Y/^����}��[��i1FJ�h�#�6�V=Wfb���<�"���e�O�ҽ�Y���s�%���o轒�z��,�=�`k�%���d��Xm� wF"�
�F�n�s;�i��9$co�,m�}GU���O����k�qI�{ؤ�_��G!���_Mi�8B3� нg�`Y��K�k��;I���������5�p+F�!N�������.k]�w�Vێ�<u��8�kVn��[�&�pĸ�0���6�˶�����X�	�bp*��"3��buzD�@�#���*�E��r�&�4��"�x
hB	�I�R� ��V+��D`�&b� W�$�o�D�R��)�;����>����rj����g�PXC��϶ғ���+}���J��>#�Cf[1<B:�9P���L-��uV;u����80��m~״ z�d����|�j+@����9R�����^^a����!EҷǌF��:*F:�ljy�d�\��xw}*:���("i���i��|U�nO0���GʌO��YȽfhT�i�1�m�a���*������&�b�	�4U���ԕ9V�=;��W����o���1�v�_6�;�u�zMX�d��p�h8T'6�a��	�����6I�,�el�Z�^���i�\-
<,o�W�=�#����1�-��
�*����㫿�s���M�2��@�٠*��)�R���cr��pt���`vd̻fßV���]�W�)rH�3 ?�c�4�����}�s������"��������)�RO&>v�� �R��q�9D�ϵ׋|��mu�D�ݰivT�j���������S]��,:ޫt���(������C����
�������Q�8����u���X)�A8Y�`��>7[��ڤ+��^�{�w�,�'BT���Î��L���E[e>��.k��6�~ސg����� �U
���`��CuT �^)q,Ӭ����5N��1�FE���u?h��3���R����\4(�b6�����#h.a�u�V[��`�瞞�0w��A���	�vg�	�{��M�PK��;�[�]'vm��Q�gj��p�X�T��I��
oٜ����7cg�&��҅8���$����ͦ��c�Q�}A�"�Å28N�ԧ.ܿ���kP�l���b �) SKh>챈Ӄ8A�.����tl��"_��="otu��=���d"aq�^�y�ǃ=Ͻ��	��ɤ�����ɉJK+ۺ�x���qx(�}��x���� ����$�(!�X����[�=hv螑̨#��f,N9;0�s����&\_~���St��2���u|��of�e��'Eb�%vEǖc�����S��ώ!��ㅨ>�b�r��u��?��w��-��C�6��S�S�>#=���hoخ>�3=
�n�7�����>�"����lM�N�)`��X��&��'�b-8��ī�f�v�D����D��N��!�7�C ���w�h�r����8���CB��o� �VH���3�ܕ_��h��ƞA��:��F�kĢ7�,��	���GZ�=>r�#��$�Z�3T{Wz�=T�#�T]J��,�O��r1h򜄱<o�P&Q��>�c:Bm+pFv�v�'���67x��y�@��`WyՉ���rA���О����Z�/$���0��.���Wx�RRC;PC6��Z���M��F4��I��-�
�#K���x�.�H�|��k�^�������b�:�ҩ���hR��I>xrj�l��,��.� 8e:��{��
��xN�A�����1�n��b�E�@��e��ݖȄf���@L��`��+���l �iSyU{L���SY�v@��o��G<��O���Ǐ8�y�p�N����x]u�����g�1��ݫ��"|�h��ز��X�Ny�=���E<j���Pb��cc,О,��g����� �[�Tj�]�Ռ3|-�c��Suu�)�^��8���I� J	��u��${M���M� �VP?�^Z�J\��է#�h
�o7�h�Ϋ�f	ʐ��*	�^�?MV�p��!���qPI��4}E�P��rd����E�(�X��4yx�V4S�.��3����pP��� �i��F���jB��)��+��y��o�؄"�=�u�|o .�z�#�x��b��+S���޹"׾M�)��m`��	*�<7���!p=f�����(y���}�#���k��Z9w��J���lU^���d�8���;VoE���.����)A��!���;��/ϕ!�L9ʺ�*'�z+{�k�"")�{0+w�w�Ǎ��HK���K
� ���/��B�JM���������snA�E�	����G��̼w��W ����o�f=���e5#)P�H�g����T���޺��⭞���"Y8P�D%��Õ�)�ȱ�w�@fڱ�5�@����f���K�;���!��֛�>?�d������0���A��ƽ�8�g���v�D�m�X�=X�Zq�8)�����*OK�/v����9�#`�+5U�4u&�U�t�8�n����2��:;��ʝ��eKõ�i���C�z�P|	� ac��Ŗ�y��8!�P���l
�pR(>�}-�4J�7T4i<*����e�vO�-���������Ix�r����0j§�*��&��t�
 H�j�׶1�fA��?l�H�x,�-e��xwɋ���U%�.�^6�&y\O,�����Ak-,�=���je`9�K�NϚC��5'�4w�g��vcu�"B7`�˞֣}b�XV�q؂�D<���9�f%���!<�(�.bІ�d�����Aq�_�ԅ��D��"�ʵ�<�w�A��$XFeB/�6$!K��\���>�.��^̸�����0�7Lw��"p�b�6u�Ϝ��[L�>u�`F���!X��a�zdZ�%��?^v<�?F��`	X,�8L.��$9�h�Ëϭ�G�`b1���
!�k�bdK��r�?C��p���'�1��kNu�+j=,��f��eޖ�T���R�\?���AEB.�렎~I�\�ʠ���H*�!G0���Ц�䈠��
1
���a��B���-kKڭ�3T6	�$����g�"ro���<���(��������F+Z�h�\X��x<�
���͉=W�����gź�H'h(�@+�6a�UGt�X��bB�X�泱7��?,P�ۅ�{z�2��1$�2��%�e��r�2D��2P�10k���Z��A� J?����A OuLa�3����"W���*�n,���y�V�b�<H"�P����b��#����#�%�ݟ 
I�|l� �;Z��O��Z�-/y�t斴���Ҷ���b�N�h�|��ݨ����v�?�k�<$+��	����i�0Ѽ4a��kJ �g#���SkDz���{ہ��=�eƄĽVGF�ӗ�H"K��"˶&=���R�M���1V�����~	@��d����P\��BA^����f�R�ٕu��\q�X�n>4&���%s�!4z�Y�����L��0,++���B�f5-�pnG6#k��,��;Ԃ����s8m\
{�SzG�+d�?�FG��ox�_Ra��!u��yӓ[J��N`H��I�$�i�n�=u@&'o����<���X���̆6�qzQ]��2='Vփ���"[�W<L�ս�r,P�ר|IxfSm�b�7����QP�b�s3� ̍O�h$x'g�#W��b��n)�(�<�s�ES$4���oÌZ��B��R���|�ɚXq�/E�Y�~��<���X��s�F��2���J���~),e˛"��ߙ����У�M�7�Y)iL���Y�s���t��r�[�L���Nw(:�&é�qu^С�;ըT��_q-���
3�Պ��jxi�I��1�%`8pw���`>ӈe�ϻj��tM���o�9�uz�PaD[z�����x�=lDǩ2�QP�B54�'�Æ�SՂ͝��������E�g�H�Sah�I$��8Wϒk.�S*�����	5��Ynt�?�Ok*�~��q�����n�N|��+%��k�!�B��v�r��u�X���"�~�� 9�y�ٞZ��?�z_���ࣶgt_h��?Ԫ�hW���w�}%�ĀFZ���V�b,���\�5dN�<��v� ~��;�R��tҼO�a�f�Ii4K�ۏ�*�І�p�<@	�H�D�������0�f� ��`\�v��y�)ntt�룙*I��r|ۻV[o�Z$��*��R�'���.s��������@��}��+�^K�T���\Ud�H�u1��;�a�����r_�G��q���z
_��q=��y�ֆ��H-��~�x�+��d���f5� ��@��>M�}��1�|���d;��9+�y
&����8�T���	t.�:eu�"b��xF��ض_�۶�-��t�-'�\ꯋ����;dƇ�GX���ᯒ���d(.YZ :�������]%�i�.� !�r��cH�a{�S��\d�*�Ms�$T4g��F���/���IJ�dl�����~)������ݽ�յ��~�m����&�Dj��Dd����J����m����w���\M�����陖Ӯjm��wʭE��d:�,ڧ˄�ԙ������ԯ��gh���|�ڃ�M?�&�/Ti�_K7��\n,�������ޱ���*�*�>��{g�9���l��Zε�nz�\�Ե+=If>���Fh�lǸ����TAX�ڻz��b�R��-ֺ�Q�h��a�l4�v.�[�z�:��g����J�����i�Ǌag�iyZ��ػUN��0Xk�7�Ԥ���F��c�j\2�$�b\�4�UU��߃�W���^<��|Ж���1y2Z�ܥ�қ(~}(A��{cZ�������'�%"ɯ�W������.Q�$v����2Z�<�����&�3U.(EQ��$=Z��D
'�1�lQU����j�
�
�/089It��6;����t-��r�����e��AI�BƩ\a�mo��j�rۂ2¸�/z���nm����3)d�J\���T�٠3:�m�"�K?Z���*���@�E[Ìa�	ŵ��T�{ҧ���Ȓ��j���5�y�2����X��`���I�e�v�h����j��'8�1}%:=8����GO7rߞ�Va��jw������؋��%�;�V �?�"U�/�끗�UX������Њ��|��zh?�Mn(�m�P��}�vo`n?3��~o$d�a���EE�X_��ܓ���I2��9�9��v8��ڤ�Qj^><��q��`AW:c�?����4��x��*}m�ִN�3S#���KB�b�$]����{� �y!
i��R%A;�P�R������5�ݟ��>up�'��k���xa ��;8H�}�i�W_}���lrN˪
3F��~�ߒS_P^��<_V�^���3v���y��W^��(���a��v0��V�=����l\o���h}Bߺ�]��R���}���7/<�"K�����)����s���J_��+��GX�F�Po�Q�.��X��4�v���$f����
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��fT�D�CԄ���ї��Dp���>JA-�P�� Q7���!mhx�����=�,K�)o�ͼ
������C�ՐG�L5�G�6p��]H��+�1\�ځ��(��w���x6�-�
H�����(�C9Qt˃��.�=p/eƷ����pHfS���9C"m4��2�N)C4�ٜ���K$}NHB+���B����#�Qy�����g#N�c��𨈀�0��:S[��|xP�?]xW+�{�@00&��d�=��qc8�iARx+�t�Ӎ=��2&n*���)�CZ��tU�^8v�Ѩx�&�<B����k`���}��^�D���K24L��
d������i���ܨ���0��YР�F�l�F������트�e����y6N��?��Y���?ꥯ�Zg��e=RE� ]dm�DWl�m:n>ȷ�L�YO�SֶB>Z�ݭ��T1'7���y�ґ'��=C��=�4�op')�I�ԅ�#�$$6$��#Gq_��3C�P՗�C&�&�Z,j�GPŎ��ca��n5�Q���<�[0�mHZ��GKc��-;��-��ۧKu�W	D;'�'���}8=���Ґ�m���gJ���)RE6���~�3�����O�>5ݧVz[�Fz_����?p�O����+;����O��I:2&�L
>[�i�ۗ��NTI'S���p���	?	�qFį�ڐ�7q9X�f�H��ˉ � �h��3%c�b�����2NЊ~N�T���C'x$M��XlxVHYEB    b3c6    25b0������0�p��~�3�(5���n&u�z0~M�#�P��۲򚻏�ŋ�����{���a���\���ڤ[~�8���9�(��r�#���sL=�'d�%�@�{DBZ��{) -A�yYS/��4R *���9�ԓ�^�F���0���hn���mz�o�+�~�����Z��.�����vJ�#i�x��۞eċ�.+Εk@X��H3U�Y�^����p�A-���YD" ?��~/���Z.eTL��HV(禊Kno�UpnҸCt�d�N����q��N{��.�N��W~j*-���<�������� ��j��@2J�@���S�K���6���$��F:��[,�;�s����$<|F=���qÑCʿ#[��YSo��%`�{"1���ǲ��T�̯fe��e�u8[)M�e�G$q��v0�St�(����BYvFa=��ߚ�N&w�!���V���&{�g���P�i�����#MU�%G/'��v�ao���G���w҉�Le��oq��ʒO��/J�'�p�qGm��@��LHdY�6��
ŵ�غ�;%q[m����C��	;��D����b��h��� .���8s[[c5D��(��q��[}�.��	y�ozA��� �}t�����eɣ�J��������-8C�<<~(%[��1�N-h�~�@�U�ɖ���������T����%�9}6���-�N����wx� ����F ���^�.Uџ�Įo��[i6h�U����mc���5���#��he�3Q8�;K�(|��(V�3 ��HS�kT��/#M'��%3��PN��}���,c�{���� 26�MQ���n~��kp,	�_N(�UT��
>v.[u���{��?��z�g\��ΤM�wDxw>F���8�2=}qe�]�3�]��)q		�&��1���i��������H��-d%��߆3��6�Xaƨ�%���I<X�f���| �P�+D}l�a�jS]���a�)��ߦk�-�m�P�)Tvד]�#�F��A��e�q���?ۻx����X� D��׭�{�R��N�1?�]0���v�2��}���RL��#��?	p���.
CU_�,0Ә1�rL݉�G+w�#$�BX)�L?�y��8�2�.�E�7� |
R�7y+�s��=��xT�3a���u�p��~c��[E���&<����ː��r�%v�*�5������.|��!$�d='p*L��eh/�G� �ek,)��}'$r���	�%�]�LC�RU�� �����`�v㌰�<n��tm�\�|$�[�׍��8�C���<~��1�{ʭ��ɱ4����p�	>�L}�E��M��ژ~P��>�k����E!����*�Z(hم�a�^�ɡ��.��\B���%P�Z��QE��AClR���8)��R��iyx�O��v	�)������8lV���XR3�p�7�^� ��O�����zD�׸�֢�c�ֲi��`&���A}D{�������ay�-�~���Y���J#gb&j����#�E�nf����ACv�O�5G�ȓp�A?�൬���e��C� �Q��u:�8)|������
2�WG�ҋ|�fu�j���2��(,��������t�����Gׁ_�"��'�2���[6~�����ڤc�cS��\S@UD�Ԫ�š�d����wMd��R�67O;�q	�L1��g�E��}�0f���=�{�֙�N�a��Ց}��/z.d�(�)���(C�TO8�ե�����8g[�&"����w��n�X^@M<�߉�����%�+�y�X$7�D\�伜��uƊ�e��r��z�r��f��W���F��|s�9����_��,Y� Q	��bm
gZ�'��KI�8��7s�4�n�s��z��Ҷ�Ϭ�am�`�b��
����ܰC�z�?��A��~��跃�66�#G;��D3�b��-����?a\
;3��"�Y�uj'Vhh�kk;�n�� .��@�t2u������.��p�"$��#o��N�Z��%/�<Y���D������'PN�����<W�yvv��!Ϫ��#�2�}���+��m
Q�ft�քbp�VM=E���#�i�#Zu���?���] ��E׻ޝ�v9J�r9=�n���ќ�j�z(�3�0/D�}����2{��ȡV�����A��Fɓ�Nv3�c�NOR��e ����݄�yc0�(�K�/�v`Ȗn�������Ə��Y�F�F����/k��K&���lcH~1�*J�����K7�FՓ$A�=�s�I������Eb��yl5����V�!j�"@���hzhXVY�մ&��r��K���4�>�����b��F�Q��-+~�Mj��$���[VM�︈6x�6�>p&b�o���G�<�>橎����~Tv4Z>���|�T)�~�_����Y�bW�=;µ���-��%�`\� �5Un�t�C�5a�����ۛ=�����(�����]�Vw�G������8CX�Ǆ��ZC��iGa񐞨}�)��-X�H�H��n�o�����˴�D폸n�ʺ�Gkϋ"u٫��4\�HF3�W�B�/X� p��F<���AǓ�*ywDgޠ-�;��A����|�W|�{�:q�������5��9k�V��N1�}��I� ���)�n��X$���ϓ$�O�5�ĉ(����j�T�M�^��`������`���`aּ������ܷ��}�8@�0:�/����U��#��$�:�&�\ôM�A1͙���6��gM�Ǯ�?[:��E��e���v������~�eo8��|��T����7�^���8���V�(����r؁F$��u$6~����q�U���=�$
o~�K+V�z�'��n������>/pBB}�oۂ��䕌=��e �s��h,�$I:�σ-�ʪV~��
|㫗��1"J��;��B�\�:�P��p9:2tl!�p#�h��;�M5���C���%�:��:�����������ӊ�E�_�ϩB�*{;��/�/��7�ԩ8q��}'��g���Ӫ�����jxe�M��`�:��@ ��u�H>�3�/K�P��>�ƎA�˜��ʿ���ȓ��'�C��$��s�Ą�̾�a��U�O�2��WޏLd�n0�C�0j����}e6
�Μ(|`�e�wU�"xn���Z��~݈.K(�E�$*�R�VH_zNz��A���{��p�-6���bfO�P���$�Y�y_q��F��VT�ʌ�^
g�
�l.Wx[�q�"�����z����viD�U�]>�,���Pu�=!�/
l下��h��RfV�U= ���hU2k�|T�;ɛ�݊jD>��Az��Z�~s1[{�D�&�����7�(��l $�$?��yߥ���Y��c["�%�Yu��}��"a�Ԛ)��9?r1ޒ���x���wTQ�c���3�/��=�QV����2��1��I��z^g�k�T�+4�����6���0�ɾ�.8&Y$6ok��)��!�!�L�v�̿�	Vs�7�-�cݾ�ȹ�K�S�˧�ߍ\�T�A{�.�+2N �J=�pR	gQR��N�ɔ�hj,�d���������5�y��hޮ���K��}��d��$"e�/�����#Y���v�
M��P�ʿC�*7(:\mw2��7��
�̞$�~�ǧ�j���蠏h������ ��u���:[�ʃ�>L*�3h[�:j�K�A��@r�A�0�{�I�7Fq;��nN解�1�qi�	1p���:�cҳ���Î������#a�y�#5p�6���#���:�.����TL�%>�6'K�)�=Wvn�����}��+R�5���p[޽���A�q�>�R��X��Ɗpc8DN����=�[	��E�a������?�0e_L�����*���t�\�C�*�R��!���rF���i�6;��qT�N�a��ԇE�G��d%�&`z3u���\�.�4��Ze���4�=|���@YԬ�E�9/����b�^��\X@�E�� �! E{��4� z[���o�׭�c+��̽���u���I���>OgQAÏ5m:_�������T��@�G�\�t�4� J�<C08Xr�������}E�Lkx�5A$��d�V7"�1�`��B9��ϥA%�4� �2�4���'�&%ـu��O���O[��j�u���A`�t����b�!D�Ѧ7D�v�P���Bq�g�����G���.N= F�;.�K��`��}��U�[X��H�g�$滕 �E�F2R��؍ذ��2>���c�w� ��� z>��j�HfB�L3�����YP�Q`���� `�2�v�^t�a��!�**�p*��?NH2&��w�wD8����&�P�!c����(��Z�L]����_wzǛ��*hk�;̒�59�>��$��]���(&�i/�	��b�jM�l�^SxM�QF�S"�3kIO4�_8���[�zP��F�����ړF
'1�*�7VKFd$@n�S�g�b���ыmtQ����@x��)�;d$P��������O�����^�V�H9�LVi����%C��xr5c������U.`,C}�9ި���g��o���ڈ���!@���hc^:W+����[�:�+VG;��(��#a�<h��da�� �̌>:>��a�6�/7�������;5�R�%�G'r��l�G���Q*"�&w� ����݇��ѩ�
�*
�itlN�}�iȁ�k�
0�6�����s��j�"sa-��L��%�Ik�PBl*;���g�E@��2'k8�̈�:q�:
*��ǳ��u�5>9U8g����i<�W@�>7�����P�E��5�Q3��Ջ�os�7%7}��#�/�~�S��=��<�뿫��me	ϢZ`j�^�b�Іb"�Q�if�[+#�n_�)���F�el����V5^?�۳ȓċt[�ϦS�oۥD,���f����M�g"At�M��QI3�mq@����s����<�Xn��^�4&��䒂BCGjN ]�|�@�^b�L0}��<̋��g��}x���j|���p0QxR�*�a��U��[R\��Rd�v�@.���^^�t�y������A9��V��ÃR��A������}=���\�ղ���ҠR9��n��1�RL��nz�p�����"�M�a�`E�s '/.h���G\(cap�M^�ϥTg\��o���%���@���c><�dj��-r�+z	P�aB� �����^ɲ��ۓZY�$}��+�4	��l���[}p�'��EQϸI%N�p��B��l憏�ay��H�/�m&^��PeŮXv@�����䄛dFE���|�d�����%hw\JLi.w%����j��u��D�[C/v/ҷ��¦^QK�-�WҚ���h�=���޿;� Kd�jKc����-�3��Ȣ��CcMS�wq�I� ��7Ջ �g�̗��	:�@&I��m���9���瞟R-�3Щ�&f&>�K�T�b=�UWb�HB�Y�K��"Nk�q9:J��xvb��E8)�@$�*�#n�Q��v�|���DH��lt�"�d*l>�?���#Z-�Y8 *�h��ꑸW)�d��;qv�s���E�z+�o��u��S^֑z32M1�8������@Vhe�M����;3h��ӣ��W��^���9�oE#q�0��+�ɫ�){j�+����^6�i�NLQ���QK�\י/�-bt� i���$?ru�l��Ү2�{��H�^bN��v����Fʍ�,uH��y�1��	��Qv�0Z�/������%~0��H���:��QnQ��2gW�·+]7��& �N��witbo���6��[9S�0e���q��42/@�p�ycߟAȆ.<<����1��::�,A�a��8����;0�ܩ}E�_}�KK2�6o����,�+[�}젔��g7_�d������\�'|�$SPm�;-=�k�[K�;��K �hfQɚ��e�b*���VDw2K�QC�����������ΨF�H[���l��a�?��`Wg%:��<#�g_9�����Ңa�=Eo�
A�#:��ꍅpb�p0pWу����jV�W�ý=� ��+3�4�PPz��K3`|h��&�'����o'Hn9~�����+4Gu�e�*d,��@�����(�?r���I�9�>=��1�B9��9�����G�#b�N��`�f!����2��N�nPM+��!k�疈p�_����}�"��+x�x�PWB�A�}��x���4�z�ߕ%wӝ2�A��*�hA�N��.�1��c�縙t�y��1�9þ�HUeL1��Z���o�[�e/=i �w�1Y��3m����[k}��f�R�h<�ǆ���ŋ�e�R�`�{��`=ud#Y���%)`�`���/�9����|�MIlJ�u=c�6�c4��?��]�7��˕,���	����*�I/ ˪��E��ҙ��~)[�I�~��j��~y�>���2��2��7�s�Ik��'�^Q�ݭX����ᴘ�7�	<�o�H��y�AY��a��f��:��5�����ѨE�4�}@��X�'=v���ݢ����$�շ��.��kx����]\�8�����B�,d������=�O5p��YR�?U���"g8g�ޜ]��0i���?�����G#S�����F��"'�ø$��> ��-�:��W᭘�!�v�8��a� �����!z�(�$�Cwjb���z@�!�0�I�Q���۰���ޘGK�FTA! �co������Z!�A��=�.J�xD\|[x\����7/��V(foىQ�[�g���� Zl�7���Խ��P�����%���ߧ�R|Hu�t"��Z��o~�ۏ4���l;m�ׇ��L��iFV�N�H{-�os_U�`���_��8�a e-(�ә���`
�[��_�9G����g��V̤�m��_r��CDhS�Z�5jJM�R�	vĩCB+F�Ӻw�@rpu;�ZE�F&A�
W� ɊPf�(��.���2����k�.3�A��������9��6���v&Y��z�y�"��5�`�F�g�խ>z��T"ߪ'�?F��?�w�O��_��A|�<v#����8�<f.��c�!����h�U6ff����	��ƴ�(ɖ�\�)Q����a�XҤ��ߋ�
rQ~�����Z�d�)����>�o�+���Aǿi��B`q���i�q#�'���Q�b���u��D��ҝKZ�_����B*�Q�ɧ��-��/�g,R���G��g1?҈f,�n�V;�Zh�#HYN��Vj����v����-�/E��#j}#{z����:��N
�w	��L���|���9\�!�7�10��Q��n	��i��Y-��"sɕ�(�[ܝC1�6�>$q�={�ugu8c7d�vd$�>7Q^G!��2Yݰ����� P�Eȕ����ƣ]z�xy��[k�S�Fҹ�h�+s<���B�&�����1"Z��QT�j���)��w������n��	%�;C	Bϻ���D��z�꣓M�J���56���v�&�����^�E�s�X1�Է���!��3�?K�f�q�Z)�i>��.��w��^b�:���9{�¸DK�i�	@J�7`�?6/�jj��<>��8]hS� 0YH��?�����}��4[��y�0p�z<5���������$%���ʴHO*�i��}$���P��(��D�"�u�ϗ���	#@a �mO6vb~2���X�+,�e~��,o5bP��l��b)��1�멙P��B����(�:[�*x�h����W�h Wyk��Ok�qhc'X�H'�8HdTH����i���Ѝ������O��Ƈ�O�ҩF�����@m��n2��Y�� \RrZ͋=^��A��cN MS�I��0�(2zyfO����6zEyjy=��Vq�����jЅAs�`�wو���%��8�z�G��5�6?��p*j���׉<$���.�Z��gu���.�9TB�j=��p*�aIu�"h���,ݲ�8~b��`F�	+�}�$��lֹTrjZ��a�n����kE��N�؃X�x6�xwX|sa��0���Hk�y���fl��?YL�獁`��.-�U+�V�|xu��	/��\M�34��Y�@��x.W҇?Y(X����`����'�R���K\gT��R�w�g�;����?V�d�e��1�L[���Q��ţaq
������R�?�����]O�&UadF?��P��]��8Ȼ��D�錷Ww��H�Ed-hM��q=��^n@K&��Ԇq��7�E+�p���.�ٓe��*�#
w'gWa�#o��[��ɷ�s.š_h�˚,Rzn��v��]�������x�4>N۠���B��f���y-"�Y3��N�؏+:^(�'>#���J� X�����E5�Ż ���%I����;w�*0n�`IX�oq�pq��IvT�@i2?D�t/�w��S�E̻���͋�����̭�X�t�J#L	E���	D�'S�V �q�Y�5"��ς#��*���	3���$%lZ� !>��&�d��s�B����Q�Ϊ�fF����t�8�X�"_oI~2�H+�\�~�f4Xx�c�R0�;�e�(����]�o�g*Q��X����&]P�m�l��C݈����JK��~�?��xIՔ��	ۈX$�����%���+#
|�����Ϙ/c����'J����`�0&�4(��ŋ�~f� D 8&��]!�`.K��)���:D��pd�xEUͼ�f*��)
��
�兓��Y�(�����-��%�א �4
�E��kn� �r��?j�����R�J[A&���8�� ~��_aۄ�a}�Y���c�҄xʪ0V��ЏV=�FO�e�PF��U�lc��R�C[���a��9~X��D��dQ@VZd�K̸%e���l0��IC�M!�����3��U��I>��vT���k��L�����]�SN� <���!�!���4�P�վ�f�Ai�T���<�yK�O~�룏�M�Cȼ������'K�p�~(��.���D�Uu>䉤�d����8U��L��I83���ɱ��"�?����3��l`��S),�XG!�U�ե��4�4Я�A��ndf)���[Z�ߣ�cv-Rxu��qĦ�}���	'�+� ��6�[�2�8�7��QxVl[��krh�螆;	X�����Z���x>�?]�R�9�]��E�Qm��4��i�������D����٠�墎p�;|?n��;��afߔЬO��h��� �%.Ê�jX"�Vݩ���8��cި
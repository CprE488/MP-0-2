XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���lƛ����2��4��!l��%��71��l��C�~���B{-��9
QcI�4s�0��clT'�>�O�v���&�e�jy0������g�O�K"�̺�p\n�B7��p�Z�+1�fu�ג�)�Q�q(�~�'��5�d{6��������ވ#�`�YP0N -�g������w�h��U<It�9�d�!򶫮��JgOl��p#��p����~;�@���$7;�r��@Xy�%���
b_d��b��}���.3����������댞Ic;�?���vˌ�=!Q�n+
�&�����.����	���.����������Ƙ�� U����	K5�A�b,�727c[y U���n�����~r"��ﬗ�Bc3�[v[a4H����e�$������[^!J�8��nԠo�0{��
��$G�]�8���U8�i�|���ْ��i	��/����gh\�ם���2
� `W��V ���ӱ�/���U�p0U۹�Zu���w���yV-5 �└~a��M�����ߪcX�ƭrM .�M���G�'�P�q˦4��p��kh�Y%KC����%_9<�l1�t�&Տ�
8�w%��4���|#=��VB6��rjsAx���k8���KװA)6����60F
b�H���.������8yd�kW��
�i�~0^]�s��o:B(�ۄ�`Ξ�ݐ�k^��}��Q�r�?��ut2$K)��c3�/":ߑ�}��I�Z�2dG������k�)|XlxVHYEB    3b09     f80�3Aa�w�/�{'��)�q�H��jD�,i�vR<�ݭ��3�r��5�]�(����������{�H.'�>pkX4�u��!z� q���-&����]�6.Vh�[P@��r���}��K���}��އ�{$����xp|9�E���1v֖�r`� ����ePV�${��aς�ʣx�Y�v��d�?
i��6{�9���X�Q+j���w$f��Z"�905�dKl��֫=?�nL}�"�M��c`��2r,���}HR�Ǯin�q�pM< n�p�U�}B�Q���1��p5w��ʸ¹�i��F^��Zt�,��A

Axb܎0��Ѓ�e�H��K=������>C��D�Ih��HX��+t7�0����æ�']�fr<�xG�hOf���9����\b�`�֮��*l���7b8TB��PL��O�C�72��<3,��t�;�O�of&n=�f#'q���������/Y����iK���!�j�#!�-b���h�C��1+��_{����g:�w�Ua뺲�>��%�4�L�SLbB�Q�6q�)��H��o-~���n�Ռ�l�T|��?������!1E���Y	g�!�Z�G�A;�?��˂;�6~���"xW*�Ae�3*�WC>?*�����> R(u� ����:m�/L70v�������٦G�)���&��;_���N]xR��Y���F/��k�8v��Zɬ{Q@Ke%��-���ţ�j$���@
��#�D<IARz�Ή��9@�o���I[��Z,��w���� CÑ�Y�9پ(�[ޥ����8Ӎ�&C�=-{�]���y���]ݪ��e��+�oV��'�;>�-]�iwM�E�Ai�-� �I���X_���K|��W9h�~o��܅�kXz�<����(,x��,���V�ql	UT~ڬ8t�-�qE�<�m�/%61�ye�¸N@n���S����/_7vB+����ȇ#m:��
̝kM�}�񕙉�e[|%x�P�P.-���K���P��e�7�8Ҍ;b�Y3t��W�x�e�o2U"���݉&�w<S('�B�q���y 3:l��2>Zb�C��U}��~A1��<�%�n�|���m�R�ڷ �����oz�d�({J���S�M�(�R>l� _Wb_�O���B��j��xk�b��y������VY=�]X�*ª���֬^��W��ݕ�a�6a��́��B3{XǶHkEntM~E����΋`?�2}��U��	pDn�O��ƙj�� ��@=�����f2������Jt����6�eX�|�co!Ŭb)~2����2�ѩ��� ��t������-״A�e�*Y<� �
o�j�7�K���2�h����`�=$E�!���S��چ��t������\���n+S�8 o��$��X����������
�)E̆�K�-dx�\��y ��~Qj��Vf���-&z8d�I�a�L`5Jｨ/X�)I�\>�6���3��
�p�qz�u��l���)��h�4�9i�s�M��k��M�Z/��kLө���)���g��;84��O���233��x$���9�L�&r0'g�l���N֊�
N�K4���KS{?Cǐ��6�$� 0��4AU�e��/�.ӹ��ߓ�M�=b��3���:bU'�`S7��&6�3�wΠdG~�|m���M L&�������Ӆ���=��G�z�|�Y��t\����"u�mUGH�-��F-Gtc��O�g�;��[2���X��i�M��E�8<� �:�
�t�8���M��a5���������: a�������%���~�R��M8��Z�s�o�/ �OI�9�f�c�s��=�js����K9>a�=e�����xö�'$�G�_ZN���k}-s˻�'#Xv�[	����uB�_H�ze7����m������-�(.D�U�]�:W�A���5�%ہ]�kaBx�]�����a��.���+H:�]�l�;�gG��΃^zZL,����ѐ	��ں�e�����:�^���l}�5^��	�d¶�={�'�M��� �ҭ���°9���	1z浨M2ڢQ)�͙��a�A���_��f�Ԝ�M��ԡ�doQt��ц� K ċ��̚��Ի�d��Ê7�s"��g��9-��x�~Y��7���l�_ܜQ�͊\aT��q��}\�6��<�e��ϋ˯ 1 ƙl]BJ�V��7��~+BMzu`N�.��ƽ0V��o��Ǣ��F�Q�:H}O+S��B��B����֝��3��`m��������K5?0��9���6?�ϡ��\�0\����Wh�v�4>e�!)��VƹZ�0,H5�8��@S�|D��C��{<�����uw^>-�	Z<Z��9�E������9��.�t���)	{��W>���󠒳�G����E��Β����~�&���r��D�
(S��,��au�i���i�|�X�=�-1H�)���S&�d����SQ%?�_y^�H$�*�a�un�*Z1}lp��a�U�p����c����ǒ���7��׏�����WLg��S� ���,lM�s���߼���`����8��65��n�p݊�{��0F\c�F�*r(K�u�K �ja^jV�]̴����76�7�Z��I�7>�Ǉ��������I4ڏM��ٝ�{y6f�#�a��K'`S�Li�W��K�]��F����2��6��YKI�K>��/��K��6�HI���pm?��g\��F���V��\�2�UOd�2H<t�5�5 ���6�En��N-2��-p��ca.AqC	!�Yv�����@2�ۢ���/ӱ�AZ*g���{�z�Qҏ$]�it(8N��]zP�-(�(6u���`�V��wC��Y�;����f*w	����a���>fP����0��@	����,Ҩ0Ôa4E��u�'���!����_mIx��#�s���~��I������%mq;�p��[���#6������m���I��I}Zc�yj���/�mn�}@�y��d��t�㷕�6�g��X��BTd=.T�I�hB^,?��U�j0ˁ�X�?�5R�)�
X؎��G7��*�Y�	A�?k$0a{���KL9���BՒ���,5�-�����<�m��Q����b {rd[�D-�@-5-�c�<�����r�4�լ:Buޫ�ЊC�:�R��¢�/ؠR@D�?�<��﶑fW�^|���Px�QH��q[���߰������	��;J8~Ug�pv���r��JK��*�C��hҷW����)���Zo���Z�<�0����A��@4�x�"�:��Bݡ]&��h����%
�4>`* ���Z��g-����0 J}fh��j�y'� TU a	��
S��H��ɽm�k�>ws��G��~`�(z�p{�\�EX����!��_Uv�J4�9�bdEm��/r6Jԩ�0),��TqM�����og޹���5ұ<#�J	�t�{Sdc:s��V}�X���,;J��d}ȵ0:0����,\�ۼΤ'h��iJ�إ2~n1k�$f��f[�E�P(�6�z�:Rx2בU�rWK�u�>��	��!�����C����%��ii���yP��)��T�Mk�^߉o�V�v�dp �}��e���S��Ϩ�;x�;��(���:����֍0�p�=.�QqA(|���%��t�\�W$�
�'������S �J���cI��*��ؖi�0�s�J���� �C�I\_7�IpM:3Y�8�="S\TLD2�w��ICݹK��6�`�'�bcz�^���#���3�9��k�0�?d5\���G,�>i��U`Ye*�"3���b_^��zW*�4�sQ��7+y
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����MB��O4o�?:��Xӳ����:��TG��?��=��5T��[��O!�Ωt�!�\M�x����ֹ#^��H�Mgؗ��F��Tc]�1Ο��~Տ��1��'����z��ߧ%4m�k�đ>3�w0���1ꌧ[^�k������D!�
��n%���!ð�
�l�|8�p5��^#����noD���*%��HY7Ƈ�����Ƃ��E��2�J��v����V.�ܵ��c����pd�<�����]L���O���dK!.�{G��d��%��4��jXI$P.�P�d�n�X��~�MA���`�c8�eo�v���^�ݜe/�D�dw�OϽF*��L������x��OO),��.�ɖ;����t۷��y�^:쒔�^G�(�k�W%�i��LhR�j����5YE�jY��9S��0@K͚��GԖΟ��P=���$���`�U3���[��T;�Tn�3"�ֻ]��%�h:��VY���C���(dm���s����"�ד<t�.����F7���eŗjx*�AJ�]��n�R�Z�G�ʱ��'������mOO"GKh�H��3�H)���4�����+T1���Ř�<��H`�8B%�ӎ{�-�(O_lw"�Ԧ���*�M�գyv2'1�|KIS�[�mv\�φ���=ݹ@,��>��'�k�m�L.(���m�ŷ�;(|�(�%�H������E��ev���ܙ��Ol%"�0N��+�E&XlxVHYEB    a037    1fe0�㭄��m��S����Vܾ4d�J�4H0P,�8F��l��ͪzl�Q���i�\���`�9gZ�H��(m(i	ʔ-b��wY��0����&�ƶqk�j �JQHPIf��^K�u��\�{k��� ���H6ݣb��ۓm�US@�y�������[Ed����@�1�ܒ���vW�(�<�Y�[�o�v#^qn�~�HN �%�/��i��_��꬜�!�ʃG����s���ݲ�p軶�!׌�yz誕0m9�gM�$�2�^��:3��&ߨ���/�	��\v�'�rp5y:��B���'���gFh�Ib�����,�Ϯ��a1F�椳�*Ϯ�Ȯٖ�%>r�/��d���pI�}�ݓ���?�(Rc��4,�+Xk�\���_G�Vadز���ˊHS>� �[v_��[�+	ǥ@`�k�YC�6�ۛ��
|�ZǲE
S�	�Vys���P���Q��xN�rM#�8�o��B$��/���-�5��ir���r3/a�d75�:m��m"�֘�f��8���CV��	�J��UG3�d�k@��+�����#�M;�0��k�	>p��SL6.(�>�S��}�8�2%zIJ�e!�5�\}�/�)��SEdS�������&��a�~D�(�N�����0��Vp'j�8�q��ͼl��"�;�9�u��	)�5��A�6�MT��WG����̙;@𱆓]�qd�ǲs�������*�p�X�u�����1Ў����C,�Qu��5o���}�R��X����v�o5!RIU}K۹�J{
b2��wr�=\�[ę��
���Đ|,F*Z�-߽�(��{b��vFz�H~�Z�+8-�
H*���TW,�Ϸ���4� ��,_kk���k9*5��m�z���:j␾�9	R�9��u@�=�N!%�*��ӗ��uW�IO|�n�A���I�Jw91m:QO��(i�Ф�Xt�
�.�C!?��|�`,.9����}d��5�X�k��Y�r�?X��_�Ū|�q�Dl+m�,߁I��J�H	ag�]{i�>�I�[.�����q"m(s�G���]�'�L�U�|1��=Л
��\6��A�Q�@]�w:��?���F���v�o~�=���-�u�=揥@|^췼��J^/j�To�?�-4ҭ�W���!���B +%��͇&�Y���W���W���O�et��ˁ�}h�n;�nپ��ڠ�m TS*�ټ�ţ����� Gq�}ZM�����
��bπL;9�}Z���̣c��xΏ�f=���%"��4�a��OW�dݠk�4M7�M|>U[���A:�VH�W4K������I�A�a� S��0T0���}�5uv(�.��y�Dc��;�,�zP�<tN+�	��G��#��&����v
��5G�i�n#���4nb��z�o�\����� ���TA�>#7�u�c�d��T�;�����H����^�]�JPH���an���*���&����68E�D��f_\���QW�Mz�0*�xL����'Z��;�h�gs2��������3?m����q�]��bY�P/�
����K۫oT&��S���8�z��ڝ����[Zl�����=�`OB �O�ݹ�����1�P]�Ё�g��bU_
�:!�H���ˁ$�6P?��q5��F�|�hL�S���/v��Qbmq�޵����y	�ɬW�v�,z��.�֚9�ӆKJ5�z��\���3�r�A��"��D�Ǿz{��G��$<������d�g�P~{��=����(���WΞ`�3����k�[�xZ�j���!2�j�QR=��O�Ա�?�>�yB���p��׬��3����8��}XX_�o�1��Z8S�i��с���cp���S����}^������(���Ũ`��N��Fvi��N���dY$�@{A=��]����>��Y����YF�3�@�鷷E��a#M�!����mj�R��W�����;�U)�v�ל��\vιl�����r�x2����Us� f�1�< }4W��:�S����j0 LkS�d���W�s��cL&]`_�gv��Y�4ŘX.��e^�F/cP�O�ݜ�e}�̮
�C���e�V�m����3�,��-S���<]���Wܪ�bÃ�#��N���-}���ds�>�T�������]�S�*S��}�x�=z������&����E�3��Om�J�v��Z4��؁X�x��&��s�,2�����+�x���lc&�~!t��|��	�I�_�Yq�P���+�wF"&���<��FV ����yLgx�n+���"���r��<=�]x2��{'��%�U˘�L���e�����j����| 3�R� ��*Ї����U���o6�c�ٹ�.�X�.��jr�C��I�~b��v�����[4�F,�$�*zZHgI2�
, ���Mϔ	DB�B�K�~����0�ҹ욜�;��qP�۹y��	γ����!}��?H.N�mY?a%�gWH_��l%�Żs���4u,���Q��%��Wjx�t�m��s�����e3�;}x�ڝn]So�֙�f�AA�t��,��1�*��7d�XhkU��p��Zb7��^J��!���*�9Ә�^�"�Rc��$r,�O|z'oUQd��A_Yڝ:�֠ğ-���I1
�����<-�hQ��c��< �>�gs�E�q�W/�6S�}n�P�2�1�f�jO�q�F�2:�df�Ryw|IC��Y��� ��H�l���3�i?��W��(T zC�l<�4�@C�5��ڧ�N�_+��l�<}{���v�R�y�T�﷿����фuw'�be�����C���98&8p�k�����\0�Z�t�W�%��p����_xg���-&L�zg˩��2��ן�� ��DS��6FJ=���W���O���
�Ǟ/s0�#�����(�aK�r�nu2�\R{5��t����t�����Z	�Ĩgz� ��������t�$N��+�Ә�ѿπ�}x-�#�TU0���2ڷ��C�qb����&�m����L/��)p��5m�I��Q~�;َp��AHJSY�~5�D��g���^� )
W��GN(��r�g~��A�s3�~���-W���&�C.�Lc�-��+}2�U��]8�?
�X�c�wڲ9�lD��c�6(���=^K�Gc���\oH^�$I��C�q'��
ե#E6��2�ˢB��(���~"dl
d�w��_w���FW��uH �w?�֮�3��-�5��L�9�]T��V`��{w�K'��1��`�� ���v����߳wOp���Ks�Y�|��M���y���RCJY��dI��-"B,ɩ����aw�'��%�Pm�X}�����[����~9����9Q�-�v�䄑(�aB��������#�թ�ds�C��$���c�����+��$�p �2/�Z.8}�or�gK�+p>đ6Bg������6E�B`&���}+� �"u���qOW��z�]��O�6��C*0y�ߜ�}��B�#����z8�jǦWCJ"��/_K1�]@���}��.3i����쏆�N!��aLs6Jl<��g
 �+%1��Z#��|ܵr�!d������۱�Ifa��H�>x$58���;�Hh&��`���u#N�����<Wnb%F�sT�8����S� �&"�6b �
�Ch��k.�f��=t����	�"��H��QY?,9Y ��d�7�b�̪��j���	�yn��C7�p��4�ef��V}�v�F�?�*��%eyW��'JcN1;�@Qش��`
�l"�M$CZ�M�����+&��;e%�����aXm������2����#�Ǧ3P�0G���������d_�'a��YB*E�l)E�͑�� |�(pA<OF&SF���v
�����),��y�����`���*��v�S_O���~��D5����Q'�����#nb D�˻�Ȍ5p 
��E^�70n7i�	�`����UF��̪^�D
2K_�uj�A/�귅�O��@���0�&i))93�~Hnߎ�Vx�:���{_ߞ/lN&�-[ֿ����\��?2;JI��4���K�!��+O�o�3�m`��^�I1lPw'JY��'�Q@W�EvP���E$��b�?�*kW����b���9P�K��=<k�5`ʫ��j<m#�w.@]���</�<�n'�� ��_R�F5Ti|0���.�82�Q�t�S�j7s�mߙ��$�;Q�Q�9`_r�k�p뒲����;9�q=��qr%$��Q��_"�GC��(�"L��Bwy�����g�&�N�bO��EId�����wGɑ�B��wh?���J��W�#�Ѣ� �����޸E0ڟ�{����8����
�	��q��:˷X�U��?��:� �,q9��`����W�ÝFs�k��c��cX����a;'�� Y]�A0� 4>���gUKD�H�m��׶^���t���#�S���B�F��/} L�Ok��wU�\���=7��<@n[�5����%����O��5]�o/;�c�F8�;�U-7������a���m7/�^!?��D�9*=]GQ׍A�����]���+��ˢ��qf\�Ҵ�(�YJ�$2�3���A�Q�`p
�B��#|Z�K�վM�/��w�ɦ�����U�4.�_�j_a��61��k�KJcu���w��o%KR:�Q���z�Py��b���sUcG"��W��>�C��:B2Hܶ�ƴ6��)D6��B]������3����4���|k����a���X@ܑ�%$/�ٳm�<��Z�0��0c��oi�G���PU�q�~�&Y��f���ed�l'8��
Z[�+ը��֣M'��p���" ���c�w��}D�S@��������Y�YI%QC+~PH#�x?�­���,���ͽq*z���dg@>�y^|?�����횣A�i���;I���u�X߷�>�B>#ΐjo��13D�c�J~�z�p�����O��":�J jn"���[=�t;��NK%؁=k��d�tt�r����s2[!Aq�1 ʄp��wnX��� �k��fN7s�����{yr�k��Ι��۠zQÇ&�e��h���C�g�;�(��5��o�z0�Q�����'��|PG��J�}�����[ h����bT`Y�$�9�`,H��z
�2e�Qff$_�6�Ŷ�\�O�r��H+ �&zC�����Ϛ/q��E�;L�-��W���P��Z~��I ��	~)�U��c��Plo�����J�pG�I7t�D3q+0�����W8I��x�适�k��?'�Jw�v6��(�����|k�2�7��g]L\E��]E͸~�i"��ؖ(J�n����s����[]�mv-t�B����S��r,��k�_L�w���ߞ�J��qh���m��{��BE�Z��z�@�D5\A�v�������a1�����1��0��a�I,4��'մz-f��M���7�0���G�Uy��(Gxb�2I�NK�8y�&�,�J��<L'ٛ`�#�4����q��a`�������8�"=, ���@2?��d�y	�\��/X"�Cf�*m�|� �۔��=Nd����v��q��.�����s��LzV7�{��ե�
}�'_U��5J�����������%�r�{�L~�(���&�:��O�\�2'>�B��:�d�k�]��°C8�-72s�I�f�[n��&�ێj9�@�I�Z XH^h>M5��
ȍ���[;u�k!	��]t����ZT�ͷ,&��$#���8{��L��Ct(����˹!Bi�/i��B��u�)��̩,�z
'�G�j-�1��ٳ���n�N�>�4� ��/	Y��n�t�hީ�c����a��C�)�eɏ����c,"q�؇�YJ�'	�x��݁�
;~~��o6Õ1��ϱ�`�83~{��+�Z������9�5a<<�����9�=I�����=��]3�\���3�
���$��g'al���㸃G�:E�-(W)&T�+����,���*N���ZN��mf:!��w��ĩkҲF)��J�Y�4&1�J�4�(��z0_[X~�P�mYĕo�Zc��W��`Գ���E`c>I%H@����R���h�)�g)�<�x(^۱�q���ͅ2@���.r�@���.ɁG<l�}9#W�x�����p_�(X�lv��l�.��2�~(S-���4kc�Ym�)=DYD1-%3�6~��p������}�G;�%�	��^�%`%���%'���[�{�!��~3Ż"��\\9
�ZG�@��i�s^ A}$'�F.[�F�&αS�TtC��.�ҡ3�E�������AU� ���Yn%�iE��o�;�=���"wB�lOj�=�pE��\���8W}^:��e1$NV���o�$h^�_�ɷ=����'�T� �����ǥm�B���1Y(�kX���#�LMb��?R��pT��$K[ۖk ��E9���$M�V�c�`H�c.޷o�x �C�N2>rF�/8�%�B�F�C�$�
����4��␆�ԉTRL���7UL���	Ó��Ì�@r��8��m.b"�x�䜻���wH�e��{��t��~yV'瓇�T�TX�`�Qe ��]�>��aRJ���k��3�����f=�W�&[����U��AՑ�b!�tz�/����uXPe��(�Kt��xH�e�ZaqK'AK_ў"���^�=t��NC~�*=`��	�b]=@����	*���*Xc�O�M'�h�=��˰� ��<�q��>�k���r���ģk���;ｰ����O�I���s�>�����ȄIIi*hB�ھ*,��կ��0���i*F��O˂��^ؕ�W�����;9���-Ӎv�K�)���G&H����gp��q_���2�Ŗܙğ���ƒ{kX�2<]�jC�BLȘ��^��J���<<�?�����%O6$�%ٗ�Nk����ax�C�/<����2�
��pfu�a���n <ԆA>= s���v�vڨT�9nQ8�׍����Z���1yhq5�)>�YW����<$�(��[�#��͜��v��Z��`�;��'�9"��� �|}��ǟ���b��z�����ն�"V�yذ�*S�,�Ēh���yv�̨24��h�m�r�����?([͏�����{�����\_�W��X���H(��H��|���6�V�nh�Yb�=�M����(�MO`W�UF�z��bH��k��:���3d>
�H�g,�M�L��\���p6.��#^��v*r2-��G�/���W#����X*Η�n�	*'���d������dW5H��?�1�``;k��	 "��0�\g��f;Ev�G�s�jZ�f���
5,��x�4�@�D�`��]� ���Q����B�`�1��z����� ���fN��<J�В�Z��-Č����Ĳ��tn�U'c�y*C8��ᭀ��b2y�By���m�xBU��# �F;�t	�Ґ����/_	>��C-�/��>V; ��L�u*�^9�����Xkd5���'�
V�Jr��I�ܿ:9�)��jk(��_�3e��{�w�m*�9���M�u�k ��4��s���N9�r�@<8�������~�9��q��̗Upr����:D�覙ݬ��� ���������l�g)U�;8U���ԫ��1|o;�-���c'�:����I$��HdY	�� 
5b����?� *@)�Y��������2�cx"�:��T�*��ݦ�=<߷9�[jY��8�N�ĵsI9,>3љ%V���|�ЛC�v� �V�ẕ~��%Ѻ�����o�b�5���S�>�B�؁��l�F:n�7�Xt�p�W��"H0V�vZ	@��U�$�!}��BE�i����P��j�$B#zN��p�F"w������ai�p�$��T�Y�WYOr��և7҈���a�	�։���>MC�g
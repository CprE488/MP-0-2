XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ue�p�)�U���	������v%��j�7��B��xr�pG`��!]�h`���%�T�������.��&ni�d�M|�f�ʀ�t���[y�u7�������.�����w*��a8��q��7;q��W�6Ȋ_5b�n=�عr9:�?zBO���հ�-��s⦽.^W?ŉ��[�(=�$�ɅH�,�&i=����7�j�p��3#-[Oh2͋c�e.oғ�̣  e4r�!;=���i��ز����.�z��ׯ3Ԣ3+�ˍ�D�d��!f���4G��織Q�U3�=e����27�:��W_]�]��2 �5��35��7ʺW�m���y�s��gM���iM�\���􋕂�e������j��L^5��.&]���S��+x�2G�D<,N�SQ�-ri�K(�.t�)XN��I�˼���C����L�D�X޶ ͌u�m/?�)���e^�l~;`���?"6Լk<���̵��؉���	ve�u��_X�`Sص��l,���1R�޳��N��&:���Q��"Z;B�J3�ZG���؜ƒ�5����6L	��fw:��+4��]��8n��RM���z��d����#C�+��7�
Z"a��X��(��{) r���<R
��O����?Q�wp.���˿"g�ܸ��.5���2�]���;P��b��'+��V�*�R�``��>�Vq*7��Q���*�&�p���O���m���r��i�j�.z��XlxVHYEB    6014    1840�>lsv��	DY���v�ϸWǝi��_��Z�R�I���T����ֳ$�-BP�^*��ET�m"$C����9WOȋ�;�cz#������M�N�m��7j��(zy�DB�R��UK?����v=~3�n��14 S�6f(%�+�;���F�RI�k+��њH����z�x~[�����)�)wu�-<UM�>B�9�u�g)���E/iQ&����Av5ia!^]|�Iw��\�m�&���L��^no}tg)H$2��7ߙߪ)#O�]��0wH"��#_���k_H&/�'�S���iE�GUM_��q~�v�K>�?}O(���]إ�l	1ױ�X�՗쫑��A���yԠk`�ꥎzh
���9��u{˥�H1�k&Y?���	�
�ᖹ�].QA��X�\z���,c��
:1���ӑ��=fq$C�.����=�ln���1/o��v� L��G]�揝X`�XMy����¼��>����4� n�����]����m�<����w�د]{���%z+"�EÊ�dx;l{-˛-�ؚj�Z����y�-dP�C����蹉d:2�XE�tp�$�b[���ؽ��z96�v�r���)!jV���2*�K��Oc���?��v��O)��-�t'���ڍ��{�|����8�PQ���.������L��Eo(��g�i�K0�r�!ґ	>��ߜ��N��{��ׄq�_W;��8:jh�Fَ:��@��9(�����R���s�ر��h>�G�f��O�=~�tYգ:���@ÛTF�u��x�}?��B���Mw;c9@ [Λ�*�D�5�s_v���L�$�U��	���i8m�Ӣ���=?;�4�^L�0q�����e����}�T�w��2pk:~䡀;֯=��ANϢ�p���[�l]�����h)�/��`���HT��n�e�����md��#o^$����e���g� � ��mj~W��9a;�K,����P��B��Z��y�~i�ZB�N���H�u�!�oUW]	g�)�Ӥ�~�\ѷ>ɗ�w��/�;��awgp����_^�׎�<����r�޴�i
޳8���~º8��{�pB���.���f���e�/�^+2��6��?Kx�\�$���1�H�)SBUT�M)]~~\��q��#{�n��y�����6�`��OA���ą�����:��!a$��Hxzh�C���˿w~cʽ�8�ki"[���ȇh���Zs��� �˵k��_����H�4"�s��^��2�1o>�!��6/�'�"���L�ھz'}v��s�.� #s&��`\3dc�/�+&3����4��w9
/Mр�3�.g--)?~@P��fy���r/Z�yD�0��gc���?�G�z
��Ļ:{�7J�u���aU�-�bg�F�\˒�@�H�ڽ��l�I��F~:�w��ڳVyM�ĦVFgih|ի�*1=9!;�*��x|w>j`��aV=>S��(���$eHm��ۘ��v��zr+�n3��wQ��8t��'Z]��	LK���t�n1�I�e�#�d��W�Ψ!o�YQ#����&�$DjLѽ�sTc�R���!i�R�/�.�����'�jW��~���x鐨�����ص��G�/H*�G�K�k���d��rE�8?,���U��D\!�n�"�
ܭ<��9�;����=��i�b�*F��˚��L��bΆ �\�d�ld����K.Oҏ��]�Va��~;V�E~��f�Ri;�K��?�����"�z���LV\a��/���>����E�-4�6����b�K����B�?�bZ��tB?�d\��̈́��"�\ymӏqf�t�>e3U�&�G,��9�����I��/����"F�us��ّ��M�U���7Cy����+z3�g��fq�k�Թ��v;�P|5���7�P�ʩ�jh�ب��1������tk��a_d@{q��6G�n<���iӟ�����]*��l��#½�4�"����J�$���!H��s�C�=;�!����s�q�1;��aeS�.z����lzjb+��c�cXqb���07�a�]t<W"v���:g;�vσ�|4Ѕ�OM۞��Wg���������:Dd������N��.�,�ɕ3��a�uS�˸�o���˙��e�p]ۄ�UM
Ǝ��1ZN[� 1v��FVn�Ŭ�N��3�&��Აr���g�"�&7�����{�E�x���N���tMq9"df��o�R�	��r#�;�L�b�a�HoR��{��E��$�]:$@�����~<��"y癢�5T�|���{0�_(��u|j�rX�N��g���Z��i�`�{I��]vDv�z�?���Do»�e�U����
��t��#l:*�-x���H�5o6���1'S�ݒ�+0�"���vO��}n����7�'B����n80�L���s]~k�{�Ӟ��Є�,>����|^�-���t�����輵2�������pO�I������O����\�.-�6�����Ĕ�����RBY:��C1y��w
U�Πfk��փ:K�+�PC��OI֕���>ӂ�����<T;S�H���CQ����<.5��4�%/��߁�wc$�Ev�P2#�%��M�l����J�����=���Mz3�J�T�)�x�q7g��Ef�1�V7�E�m�_��2d�Љ���1\_J��Dƅ�?��}�̉F�w��+�f���`�>Q�:�Ԅg�r+�TI�*�8͜�z�j�k���^s�^e?�qB��tU�
7
	����a���n�/�c�4��=�
U������o0/�UY���<�]9��|
Y�'���7i$I'&�!$U�_r�Q'֕�2�d��vu�N�E����:��5Y(î��H�UjAr���Q+��o������=ƈ��l��CF�k�=�w1�5�A�A C���HS5d�|�q�.z���L�2ِD�������g��쒕('���/��Ͷ���ǻY !P�J�pl)8JkU����P 0�qd�Y��0��V��A��Q|=g@o,�C�������M
�5�ji�W��۩D�<ԗGSCqkb,���*��#z��7E;d�۟�����B�6%����۬�~W�*{^'(��o�rZ�c P��a쌀�a���?������.�K)S7�����^�;Vm�tB4[�0���κ�?ӫ93������.�^��Ma�A-q��=�I�s5�ؽ{�0���$������=���'�ZB.Y<�/��-o����_2hZ$�J���V��v{�[tڵ3���ph\P�3r���F�<(����} �|�]��v{�6��]�1j��89@ ��p�jX���^N���R`��_^,�`>���͡9��X�Ƶ6����l��?���_���9��>���3<�(ݷg
F9���p.Ri?H�z�^ĵ����O���x��T�)���e����NL�:�6��vP��b�I[�]P�1�[��D���>Wn��(�ğ�OL9�tח�.ޟ���_�Q5�b�̌��!;L�����C���5t�\�?=��G��ѵP��s���g�l	cM�b���)z�,�p�s���7Ƹ�5�����Ԑ�y2��R�΢�N��AV�����Bõ�o�\�)("�q��� ٖg'>M,�*��,�W��`�֖*-���W���Ǆ[7�satz5�3aH��^۞^��4R�!���@��?~UfA�KM[�w�cI�3�� 8r��X�f�;�~Q���"�p�+��M�M����{`�F��bs&�mm��J���z�O$٩��{��b����Ϋ���RW�r��6�������<B2��8��M5�w�,!M(@�R��s�Hu1��W8r��ҷ���6�X&&h\�4Nf��3��#���Q�A�<��l���Ѿ�j:?v���$7�W^�C����o�ݧu���ŗ���dxm�B4�@���V핏
ΐ���!�3l-I�O�n�J��3�j��쳋��3����}�)�ݛ��?�������6(ul+�ў�p�� �1=c���|��z�oI,1�#�&{4�z�>/�ԽoY�Oh�ߙ��F��l��������7��Լ6��1G�	0 �r"_�	R���-uA�)��+&�x���b��Ϭ�C��'?F����R{\U�f��4߀�U�SY�o�)��d�����M*0��Nds�{ߒ�f�4���aw}Vʘ�a���`7�e�@J�Y2Q]1�*���	�`��h0�3�1j�G��O����}���j	'/sB����׏��ȁ�+=^�n+�M��Ǣ���Y�����Q�3�[0�{�u�o}?��|ՆCRɟ���Q�Q�9<�6(�H �b@I��|�LN���,M�Oa3�pE��e@}[� g�q=o
b
���owq�w�:���s&'?9i�l^���]��F�!����[!���dx:N�ɦS�v��.���x�C��T�K[���}��P觐�VrgD&l�B&*�̰��� $������?nd���*n�#Nv��C�ڙ�jA����TC�3#!�R���5�j���Dg��C;��kR�g��uFK���\����[^�Ec�W��_X��%R�M;�R��6�mR�����<0��&���.1 6(���8R',X���ƽ��VG�1�&��D�t�B��ɿ��J0�ڟf`,]jr�u�r���_!K
���"ȩs�y(`y���La�2�~8������gS�W�!#���P�s;	),��+Cj=o�$�}`aK�̮�U�1��Z�C����r7��.i������88��,t�R�J��:�{�/c!����+{���$<��An��cx��@~���0�=eOZ�NG��M�8w�]P�̠W���?@q���T?�ѩV�H}�m*˻D�m�}���D���B�b�)�J�F�2 ⠣~������/������n�%���r9��F�\�Āht1�_��k�%��/�a$�T8���oN�Tr�w��<����s�x�"�a+B�&�x���|T�ӡH��&��ˣ����e�<�3>t`�*xg�4�����$O�yOc��8�ɳ�N�L)��3�Dl�ot��d�֥ᢈc�r�z�+�F�K�;�i�N������[��X�d�L�P.�l<{U#:R��h�8��yh�%m�pX��OmKI�x�Ԩ�]�n)���س��:���(ȗb�<���{�$�r!������%_N���;#w��bAJ��"�C��)��[�<��ٗ:Ej���⓮�F<�ޕL��]�p8,w2�?8��i#�[��h�G�Ut<�m��!d&p�e(!:�2xn|B��=$���@.?'�`���>����|�Cob��u[7Q9��G �&)�2��+��`3:��`�*/���2<	��;�kS
����2���|�0��B�UjL�-�{���sQ�a��/h����6-~3v|�0`>�m�?�Y�/�C�κm�ت�,e�pg8���m��+/ۣ�I�
��ר���� *��+����[~����G\�)���?�����M����%�/)�� ܓs�k�
U�v�v���QWx򒭢.���Ϊr�a�k��`A˗��|��z�N7(��e0��]Z>�w�䣿�yCG�!�0��2ԡG�~\_�"��D#�� �ekL�8u��A�٨��̉�?��J� ]����(�q�x����Dl(�A����^�c�<!Ʈ��_��T��F`'q��n	��Uj�'e#��Sm�g��E'�[U���(�{�����a��׿�,�F�)�V��%�(נW���>_$��	�sp%���/��n,���a_����p�5'0fdʉxŢJT���#�b�@����w��8U��ѓ�r�=}��].r����"^�)��Kl\큩Ui�ԍ�;��V�-�Ďd*@3�'3�پE>=���^ʨ���QzA����
XP����B���8~��AZ��02�Q8��w��'�9ծ;��bfG��B>-F��@��J��J���^�z��@�y+H��8��	��r�²�u��	�&��v_��Ia����nr���9��5of�gR�_"�9���v�;��"���:){wX�K~~�
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0��0�q�[�o�`_j�J9�ha3��-����]�d�p����-om7NZ��&�[Y�X�~1��Y��ia\E0������I}��y�Q�w]��������%W))��ױI���r���A�ǅ�-�/(�Ŀ�x;J�Y-���X�M߱��ގ��\�C��-K��w�@/��{��-_qB��/�L�{9��7ܦ+�r��9�TN��Q�]��_�#
�H���l�ෆ@���8�9���0 ��6P_N��djT��*�*�_{�ian6��^#�z3��YTRhkt<aB�*,&�m���*�-8k}K���;#��m*Z#D���*�H`����u*�m�� � -�ذ
xc����y�������� �{�vRn���]ܚ��}J�G_�N7ZP@�����_ys/5₤�N��ם��lvI�2�b���ס����(���
��D;[�oC���Q���'��ڶ�|wou[h;g�/#�r5�E���Gљ��N%���a������Q[l$8l%��݂�'͔jy�B1�������_B^��O��k2>F��C�W���5��&6�O#��?��] 0v��l#q  �������X��V�>^���DGcB�Av0��O9�*vӪ��V�,�9*�yy��S��(Zp��������wq�kV��<����W[[1��r"�d8�6S���mE2;���$�a�i(�����	�n�x�P+*-"\�Sjbլ<e���9�!��t�wY��'���j3��Ăw�XlxVHYEB    42ae    1110�kǖ~���\��%�~ g�:z�h܄Ö�=վ1����(���`��WV�����ЈV���rU�-,U�K�F� ً�G��{��e��ph��֔s�*�J��葙�F|�M�����ZTl[7?q���C����=�z�����&TÔ���G��l�[�o���CVa��z�PxT��S��w�Xo��a3K�`�T���q'���
�K�;oj��H��S�z��b��#�NF$���*���X�v��eO��|�,�*��$qJҁQO#�&���"b*׼����t�%/�����\�k��*����s 7�l�V~�@9: ���	ʉ�0�3Z<!6��O��eN�A]���㞦Zͫm������0��N;4�V��s�4�n��Mד3��W�݃>��������X��?z	'N�\��n�D�����P���p�ýZۗ�j�i�se�&�r}����6�����P�U�߮ЏO[3�2euq�bD�������˻��� �fS,��x����a&�\�M�d1���;D��L� �"".���ca�{,MG/�&�����aZY/��2����Y"�~>�kiv_�i߸0�l��]��<�`��v�N�}L���8��k/d�Wt�X��	g������:nn᪭���ʛ���Y���1��_�����[(����R���i�'�g}�5�����eb{H�|�ƭF'e��!�h�{f��~}B��r�sd3��Y�MŔe��YWwNW��c�l��OF�Dڅ�y�V"L�ƧT�l׺JJG�=��s�:qsd?Ƶ�qN�b0׾����5�|Ic��#�O��l���A�?Te�ۃ<����-K�C��R�,�'C���j���q��5��{�E�"��$�K �(��Z�;� �w�vO��\�Ձ-��c�����f�*�bD^6qJ�7Ow<��u���Ө��7{D�P�u(��u��v��E��4-�}�@��5M���Y�q��`d9�㝏@"��a�J�,�*��;����H����l���U�e~���}�����U *��qs\<< ��_p���i�Õe��iC�C�}��k�x��C}4�lYz�iԀs�G�t���q�џC\&�9��`V�&��}���c5��<wi�OhqF5�����W��K΅�+��u%18�L0�f_q�=�0�5f�pi_�i��U?���޵�M?Y6��A#N���lg���gN�������/p�R5$�^�o/��8U��^`6�
7�{�UZ�®�Zв����r�0/��6s6i��Ǒ��G��(;��Xc%�Ի�ﺩ�YT�����*K��<��eA4���	<�k��l��X�a��qa�j��zR��gQ��[BI�	�?�K��Q��و�Qv������~�{vˆ:��F
�a��)�&i��K �� c�$��e"F�O��r>q�Dؕg�R�R���ۮ� �u��1��}��+�\Y,+�7*��P߹�h��D��g���8z������p#؃�nw�P�@;�"=�/_�uM�� ������V�}6�����B��g򬵢��e)x�P���!s�Wz�K���m��3�چUN`��������XhFP2�����6�c9ƺ���$Lմ�S�e��4�8d՚S�<
p쒮�d�δ�a�c>�T.C��k��c$`���6��5�#��
=3�2y���bHL0��6E�u��m%X<2t������W:2��H���ǘ�Q��`�$�����[���SP�l~Ot)�>��EĈj"�1ґ����vqv�����Г .�CV;���U�+844�ǪӼ��r��s�y�<{]�5�U�����2t[c���r����H��Õ���a2�A+�*��:�/y�Y�Z7�����*�`���Q�I2�f ��V�nH�g�p�L����7�S��7���
��#ڪ&T&���Zv��)b�V����WJ�t��b��Z�a��N2��
'��n*�s��i��g<��`����&��\W���
׶q�@+5��;����
�Gl	cV_q;��X���̴�%���|�:εPP=��\|4�Ţ�r�þ �(� ��H��k���\�[%"���&�_>����CA�����0�8�+_M��Q�@�\5��76�K�oNSq�m�G��P�&t2V����K��ZQ'=��$:���=
�8Δ/��q�j
�-��kD�6 ���`1fa��$�}�fo[1%R!� 僯Q�!�;�!�&�Gc��]0�#~�3�IN��X���!H r�g_�c��N�
zƌ��I��J�/ Pc{e��X6���m�%���P�8�
�S���cnoSP����vQZ?Y��$f�*�t���8�`%>%�8Vͷ�j��o��L���W�UOe�+>9D�p)�E��%���KdA�o�hb]W��݆�GL�bz��S@	n������$��i��F��[��y���ꝫr�s.��%>^*L��l?����ϼ��[d�QP4���m�!��ߎ�$�ͦ��/4�tx~' ��>!�`�0���;"������+�a�,N��v��ǻ!"�Fv��d\]*8�+M@�ZdY����k_�?��Й� �E��w�	�����yb�՝0+e։��Ǩ �N��R�:~����4 ����_��ש�`�N�]�k������w�9�dcg�Ѿ7���9yQ��>���@zK=�P���F�ϡD[6.�$�9'�_+���u`����m���&n��wPLo$�����k�"����d�˓6��e)���3�B{�J_�������g�T��J ]E��b9o��7�
@O�߱z�|��ʋ�	]�n�zm��f}�_�7����\�O�p�Z~i�b�S��S�t�p�V2�P�@�fx��,T�v��B����Z�=���_ �]��I�;� �t�B_ ~�y��.4� ,��2�a,i{XA�A(��y,"�FGF��4���YEZ]?qp(!�Gh�+��������&��t���{��4�����d�Y �q%�(�|g7��|읥ڴ�|��ꋰ��ތR9`���[�#^n�^�ㄅ0�[*�j��y",���ݺ�?�z�	�32b�nAH*����/ ;���	��������k�$s�M��ݚ0H��X��R�����]c�^�l��l��� F�t=�<������U?��Z�f�l^9T�˴�����Oe���^l����3ʧ��L�z��W�mX+�pw9��>g�<o��gX��0�%�!��{��:�t�~���z��� Wl��R#ȏ��f���/�B����gܿG>��:�:*���6���mFq�$���h�X� ��Ϟy���zL�i����'l-%��:��H��Q�� ����E�o�xf'��9LCҏ�li�8]�>}�Y�HO�^Y�}uVmCsr�+F"ьMN/0�H���l�%70;pK����=v�,t��\Fc��(:�^];i')@	��
��gZ��us�V�7���Mu��Bz�����İ��>�x��!L=��C?~zw�|#^ܻ`�����I�q�!SMǭ�Do�(p^��>��!|�A��S�8���vr�=�ɲ�Y|O�}��)���`�c-H�u|!�1�Ld�}E�>��vYF��~Y5A�����=I�m����kkB��5�}j<�V��-�X8�� �k�Pà8DB���c̕�}� ��Dz�*M����n�!��Z�ͣ�ؘ�����M0x��i}�*T��q�!��cͳ\8���1�ɧ���L���:�:�| �a駕���C��v������/�@��҇S>S�Q�H�r(��u9�^s�s�O��Q�3%!t�Ny��}�欓�χ��W�4'�D�ʘ��Jt{F�F�q�n7t	皅�1n!����oq�1��}# ���,�];u �����L@^�ZT,��Ƌ��k�GEi� ���� =� P���s����D3 o�4ѠX�oV�ɝ��l���In�y  ;UZ �`}m�����K�*��U�D�'�"*2{=J�f���n�#H�匌y���P�'�Z���,t��^����V~P�������t�8�kꃋ����$ݽd|]�ˡ�;��Ֆ��~|E��|��S��C�2���~SkL�YP	�&#���E
�c/����8��N���OXg�3�j�_Lc�Flz�
K5Ȭw+�f"u��Q4|��<?��7K#E5!"`.�KPh���������[�����ߍh�n{V8K���ΪP��/���ٵ��`>�ۋR�ދ$�7�;�
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o{�i��ߘ����)��x�o���^!��}z<��u��򖢒�>�p��0}���$�g�m�Sa#�Vt}�q,����	������!�M��b��^��*�ރ9}�o�p=��p=�
��r��*ZCm?%�	+ �2�#g)Ү`LC�B�8��G�2�>���a���wЎ�%w�WCV[�0� �DX
1Er%�}�0��&r�&%�)�x`�[w�
�G��t^��X��s����{�3�c!,Y1�ы鉍�on�/�z8��^����v�R�Gr̦<^�0q���Swy���mΰAɔV`oȓ]j��-U�m��	����x����*U^ot��_,^�^���w<
�lP�Dm��l#_���a�����!��D���N�'�����J�$"��y-��]�&��+}PcS9��l��O�ے�й�!(�?9?��8m�x~�.��Ŵ���	��6�β��r\��(�Cm��t�%����#G��Cq,^��7�Ҡ@�ɐ��TC���<w9Oz��ޮ��gJR��>|����ᶰd��|~��q��I��2�E5�D�y�-vBU��I���*���;[c�:�?�ǽ��5ϑ��jC@��^!����2������|^��z0|P���ȭ�&�Q�3�������ry�C=��Pf�[Kq���̚���֎����-x����-`w~�i�7l��T]=��l�RuG֥?����. tV��^,��;�Fl�8�#9���Vg]XlxVHYEB    6346    1790h�7j�@T�=*�Wʃ���ڻºx}S#F�`��u�S�e)]��,�������W�ҵ���4Mw�s{�'��
�}P,�-z�;F���c�Շ;Ek��]X5n��g<[3]�	"Xi	EUB3T�Bx?����KKo�
m�������@^+vQq�1��1I�he�G����,<��[p�lC��0���0 �G�]� ��j���ͫ`����Y�&JD	�i+��M>�F�L����2��;��J'cU��?&�pO�a�N�O���3���RGK󌯮v�s��h���'/݂�W��Y
�Pʋ��M5v/'��C_�}����fr0<*�? y�W�#����Ua�jV�l�K6�1;���k
�^�k��>&�Mx�'/�a����-*;���u��
�yܡ1\��>���;y������V|������8����J�fko�IM���b�<��~X%^�r-��'��;/4`u$���+���$�I,G����Ā��#��&�e��")������c�O��.�3�E�P���N��@��*�\kE�>����=^y����06��_�	�n�9��zi�vW�W��!@�Vi#���a\\l,T��/�P�qo��(b�0 ���Q�2vl�o�аN����c��$���x�g��R�\����I���j,#�s��ĴW'�B��Z ����3&�fvo��z:3+	�h�֯���)Ohb�5=D�r�B\q~��'.{03�Ȼ���t�驴����#�Ζ��a$5h��ξ|��KY�1:��u�!�;��b�WJ�?�ʴ�>c]���;Zy��A���E�%)|94�r��w�}lS���?x�5� *�����Sm���>�0F/:>1�R�����)��a�쟎��~�n��	�t�Z	{ṽ@5��rIft��²WY[˲��ëI���~����~Im%�9�Ѹ����p2`�G		�%���5B�؉T4��t�������$~x��.]H�2FCi<m3�p�I޼º����Ʃ0�f\VH �3w�����)������F��)wj
��v1�/LL�[^��!m@n}�.��A����5ؤ�+1k��7֤'��S�;�$P�
��?QLn���4�ϝ?q0��r�1;�����d׵��2`�7bi��F���2���ƁQ�б��1��� ��~�#t��w �%���xw�I�y//��c��K�C,�C�_U���6�ʼ��t�l�X	<5���Y�{-rb�D��#>$U��­C0��l� `��;�6L���V����tD���R���K�ol�ݝ{;KOg��<�S-�6��Y��f���A쾼���Ɓײ���U]fq�&�ي%�Q�M���\���9�$���bU}a��;�Oh��$$�~���q�)���K�G���I.���O����?���(n�����Y�� ���:���,����睁Rl�8�_%�%��i��9�<�Xi͟p��ub�%�E�V:�kS\߫����ہ�*s�I�_̈́ܕ�?�$/)%Th�����Iӽ#�%t�gC��oB�=$��3�j����v�����-�~)~�仩�@��"j2�3ڮ���}�ߕ�l ]:�
4]~	�H��A��md�9�����-�Z�������P+��Q�
J��s�(�;ԡ�h��!��fU�?�ȕ-X��RqJ�$�8o�I�,+�/O�BZ��o�
Kq�r�~�����ˣ�������dmJ�(4LX�K65�7�o������U�(�r:���k�8�)�c���6�UڥxD�I��iG��}�@c�a��J��2�!臵3��x8�.�����s'T02'�;�j�� u�g֞�u*�s��4�T��H��e}C��s���N@�/�THJKs'Oٸ��ddx�|��������P�1�!џ���R[��+�>�ٞ����f���3���s�?5��1Ʒ�Q��a!9t���%Ii)-��AJ�O�!lhk�(��� ��c���j[�e���c�4$�%��U|���������l��|�{&�ޔ��&��8K`�&�,�n�i}7T���.�s��X$T�v��vbi�Cq����P��֙����bY�}^�'�K�Pb�ӳ�!<�����lK�B��}��G =��:�_���D�qX�EdP���g��8��2 ���&F�������U,R<���P���jsl��9�ս,�{���"��n����U����"庛�0�~A���aS}�0�i�O�v�����x\�e�PS:�cOM��>ZW��t%�����&T���.��N1V�P;��a+��?oB�o�Ud��E��J�a�z��
M*�ȍ���!� L@K��_���k�,�,-N��4B+��,��+H�^�����t�Ԁ�/
��sy,|�+��}�0�u+*1�8�(�ģj��PFy$�����e{<��j๸�@)�w����E��*�{�3}�c��!�2������� �ﻧ���_t�����s��b2�F@SL����N��V�{��*��|������q��Kǻ����i��t>�&�h/_KSf-�K��u	Z9��m��۳٬mf����ـ�O�A�����\[�ڿ��>�e��o ��]_��ćυ��z��,-�l������y�5���wnԦ����7��W3tB�Eh�1��<��0���\�d��}�Ќ�oX�n�d�I/��P�q��\�'v*e<��MD�9w��?�L�NEBv���	9��~��w s��Aǵ��m
(��m;�A�����"$���vO:$~q�' g狒��I{za�f���=���Jj��ަ�^�j$���;#_�A����0
�j7v{B>ܘp�&8g��[��3��t�62�`̐�i��E kC!=� 
(�M��:�-W����Ҿ������kXs>��uԠ��j�A�L��!M���`��Xv�l��O��5\W����jPk��qH3����=hd���j��2���f�'&g�I%�^{���3�˗�	�R��VBid�( � b��p�k� �S%��zq}�!�[���])�eP��&�G�8>藻k��=�,�x�I�JL��L@WYT���H_� ����A5�����%�`#pUV�1�J�r�J^��1^��Y�Nu�$��K�ؑ��M�`�)t��q��_A1���{[��=�Ɂ���:�,���aI�K!EdS�(TAc��4��c_
���s�>�cqt����.��_<�������	�S*pE�:'�4�����[G/ysa^(��G`ZAQ1#��
�6hwׅ��꾼C��B������)ۦ��7a5��B5���T�ħ��2�&��E ��~��ū-}L6)/H����s�h1z�>�$����j`Ȩ�i�w꒹�'���m��HG�{}�M�Gs'M���Q���Ǐ�W��Nx�dOD���K��c�����������L��N��dԮ�W^Nj��%���Yy�d
�ޙ<��81�!��c���e��x�y'BMq(/b�����dX�"�*-�#)���m�H�{⤖�G��o3�ig�?b��j|z�@�,�4�Ňw�E%D�V�ó/��>��&ٕ������P'�f�O��I�Q�	���&��{��h$;W��p��:�����Q%��n�� ���"6�<6+v"T��Aѓ�N�H84�eF����VO�,,@=3�g������X*�t���Q�w���b�����7D��D�k���+i!~��y��u��\a�V7�ԧC�;���nm�<��E�F��YUP�
��,�^MLI���V���r?�L��~�7.���]T�+v��m�=�1���q�M��gH��[�y}�/t��$��ɺK�v�Ez:lqr0ɄM��|[���h��*q�Ͷ��1O�
�I9D`B���}��~ˇ��h��/;Ǽ�c	�y������v�4��Q�Tq{z�=j��ێ���(J�qv)�L���q���Z���9/���
�k�b�c����#�}1�ئ�U���6�����8����>�cO�7�(��~G���H����j��� HӔ�g������&=ŌZBm��};-'I.��;�6�^E�ҍ[��o��^ܬ:�6�����u�~�_�o����hhgY$����pQz~^3m/��Z��ւ�j�~���ƚz?�z,��Z��*�$n4�Y7��,���qw̬*��as`����R:E�]�)�D�3��J\�f�n\�����^��Nh�������T�)ď1(6k�wR�W��S�k~&�<�gf�m�;���݀�'J��O0�i(����
'n+n��n�K|�3��#�r�_�zmc��0m(Ѳ����fAⷧ���8��n��m@Wa��.iv�suV��}�:Z��5vm{��}gZ��z���qѪÅ����̈́o�ܣ$
I7AZL��Vp!F�L�q��x)��m��~_�IpBHv� ��q��&f�~����$y~]C��`;c��0��A���r�O�F���[�G���� �JK3��w��-ﴛڳ\����
cz���1d���Jcn����P�gkK�|�d���YՋom��I�kx�Nj!���{�J��U�?&!ha�a�TGN�b@��|��!�go}��<�j�� ֶ7��"S��?��o=��\�{6���"��ԙk�fo|᧵5��)�`��$�暽��.��E��e�zm�+�6/��#p�M�e^���(��ǳ�v��+s.��.�9�52�v�!��!g5PB��Y2�����r��v����N1��9PH��.�⢷7�G��o�tU�b�e�|�hku�������2�@�s�;_o�`�#�N��A����Ws�Ims�+���ùl����~�1�Ah�B<��k�is��T��r�l��o?}�"�߂i��A�k/a|�M	���Ja1H����
���$ �%��OZ�*&���8(b�hÇ`�'���a �'�W���xI�4zt�!�GW	��k�De�@F�^�m�}W�+q�B`�5�/��6���j�ǁ�"HK}�:dHKӍ�>J͔�]�F]Iv�Hƌ*N�[�G6[���z�n�r���-�
�C��N�=�ς��_4[�~�e"@���aBP�ʸd�g4h@��L�ѩ��&�Wa<��d	�<�R.'��l��;>Gt�4ɮ���W�9��ƾTd{h6>��""$'yɅ&��i�$��������U���p���㩸ʼ�z�[5�Oڀ[����ں���@W=B0�ì�Ǵ���\~~D��u%~�P�#�i��i�߼�r���Ϭ�؎���@�_g���V����sv<2��T���y�X���ָ-?h�*���f���+������I9*b�s`�G�����-���1��l6�l��� P�-�������y[��� =����^����<ȝ<�oo%���v��؏����?�w�n����풤|�^�6l�5�{�+�̢��ß*�z��f�޿�}��g7m��^bD���1_tA��OP�ÓH���F��(G�\}�r��K�����|�nK%\��J�c�p
p��! Gp�� %[�'���uw�c!�.n��_�a��Zq�
��.X��)lf%\Z\w� ���U֓%�!�\�چܖM�2 Y�f.�ǭq��v�Ԙ�Ѭ.��E\�N1��6TD�)��ㅵgs@����=.�#���[���B��_bE�o*m� ���c�*m9�'½���^�(j�z�!��c���_�Lƛ�1� ��̯�k	bxu�Pvu#jWn���-�X��U�Q5����b��sv�mPSW��Ky- �(�P!&v�]�s�S��ݴ�0�Ю��un�Oߜޖ���b�4-����pb*O��$HB�I䋃̊�B����c�u->Bח,��
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����c[�py���N�n���t	�=j�R���⡹v����pH���َ�7��a�����&=)_�h31�����Z����M�����`�<��j�
0�E��@�	�8��q��i�Ԑ\���u�i^.��ބ���K+�eK��f�h|n2A�[][u�3���+r�ԧW�(�|�p䱵ر��N�묏��2t��cj�����d��/�ot`w��2�Q�����c6��(r���Nh}B�b�E�Vؾ�נا�'v������Z�[j����gl��$����f��Lu-�?�v��0
����o)���4�}�_�`/��������"O������"!ۮ���OR�-���g҄�nL~��;HY �	�����3>�����L7e(���o@%�W�3a�Ft!�kS�%��?n�E8�K��7U��U�u?��A>-�lx��~h\fe(*&1<菸�����R���.��t	�m��z��|*�5�@Z!���^��N�e�ج��V��E��f,�(�D�K;	u'�af�sZ��d=7�؎Bmd�G0�J!���p�z�LE�A!?�{~�)4�?����)���A
d}\r�H�+���7��{�$��e��銔�`��#Au�*O���Nm�f�ˁ9�3��l�\���{k[q
-,�CIh 涿�NFտ��e�`�%��j�)�Kaa��V��m�#.K�կ��2u��`�Vj�dtǟm�rOΉ "F$R �e^���RgT�Q�}����OL��\��XlxVHYEB    95d3    18d0�ހ�ʥ�3�^�]�Q�������'y��2�.�6�B��N���[��F$vM��t�8��t_�"�6�K��8�)��Ԍ�pM���"�������)����r���U4��� ���:��[��9~h��G��s*�~���;&kw�+G[����Q�6�1�y���DPT�I#�M|º��PM��R����(7
�f�]6_^f,��.�ES�����rS�K��+U��
Fom� fô�G�0Jo}�-��ZV��}*�2�ke	 ��`�*���hz�3��y�D��S
�K�H,�[��U�<�F9N]8� ��r�()�=�[{FL�6JHd���<����h@h��b�޶�;ه؂�oG^s��J�7[�s����E�av,���E��Ӳ�=���m�lT����:�ǿRQ��7��s�X��o|˥���$iG�na(�����Ċ�T�|Q�cӍ[��m���A�0�Od#��~L�:�|���n��������(�%x]iҏ���X�r�/�(�+�)j}�zr������?��Ɔ���b��J�4����+k�D;�d�"����7ݙ�	 O����H����m	�x�B�i�ߚ��X�.��1��v���б�=i�]~���,������,��FJ�NgⒷ8�|~�&b�
r(��͙�F��_n��0Ϙs��`���Vk�r� ���}�	:[v"GR��������={HAb��D$C.��Ӫ���
'��PV~J��*WƼ�g�l��W���kkE� ����u�������ciP���WȗrS��
�0Ί~2/&o&�?�@�,�@g.v����N�b��e� T�	M�UE�{ݼ�9�����&�>��7�W��&4���w|��?��gG���n߀'�&�l&���sg�q���]�{d�~ϴ�K�̈́Q���������@��Sh�:wV������s���w�Q�)Y�E/�N�Gκ֍s��.煿"~���tEO���Y�,l��v2Fo��xH$n@����5%���	}�\RÖ���2=a's�� �.|
X+Zu�G��XJ��j������O����Փv��Õ�H��2!��8�~�Z�`D��w]�4�׸I)�tL0`�?��Q:�Y�zxw��@P�yl�,�;�#ܧ�:/ΆU�b�*��
�E�߻ٔ�S]��_�^�{�SG�93��=T;Y�_�~ �[��r #MV���8�@z=e
��ñ��:0\^X+�@��;q����]`��_��'�j�o�1h��rrx~Q�t��go��K�Q��e�]�	�Ho�HՔ_ >kwH~�W����$����E�(�Õ��DQ(��U���>7V�F,�j%E	T0\B�f��f��r�=U�w����[ʘ��U���a�ѳ,���n�
�C@�!�a���P���2��L��������*Z�(��&j�M�d-����/W��%װW��vE��4/qy�\#�`Aݓ}���K�>�,�n9�ua6"�m��"ZKnw��.����x̤��Q�0�:�e|��ɵJ��g�ω[�^�:0d�o_����A����	9�js�p�j��;��﷽���3�<�z?g�G�yz.fO�l���x)�H'�0=#��z����ñ������a��yM�O*��Bk�㻓Ζ~�-�G�Y���'�t�)�]���s�"	~M�H�����?Qf�:�]�	{�k���"ɬ*�^I�#5���J�g��4�y���yQ�y���_��Q�H���4(�3��������8M��x��T��N�GYn�Ox��w҈������U8C�R��ўųx�7�yj.x�0��x��s`Q�7�a�i
�g�}�s�H�>�1m#u�%���ƴ�R�(��"ݲ���F���}@[P1��q%���!h�+�:���md�B.b<��ս��&��Yr�^����f2$��l�s�\ǀ�,�Z��ؕ�9���p]�)�wNX*�{�9��I2�+9-�*[KPV�#�7�PG>���/|�����������d@G��ᯚ\ű`$\@@o�l��x�T�L���
�3�#��E-�{a�ȧ�wK6#�+C~��c���:�ˈ=RyRe��	̐bǾ��w5������3���tkM;~���a^f��+'S�т��L8��9!��]�����*eBE9�
p��x��N�e���aWs�c��'{q��J��I�i|xQ{kг��)S�Ԑ��K���ڌ'pG�����^�>˖EA������]�!�3tAB
��jMB�7aғ�ۼ�]����Wc�K��:7����g��3�Mx۷�r�oc�^:W��f#f���Lc�7�`�Ւ��tP�w�1+!6[&�F�@�n�����%���8 w�a�r�KZb�-9�;��t�p3j�>�7�Mr�U$#lBK;��/q��pZu�Up��]�=���щ���a ~�̔{J�}"2)�����%~�t�>�Ss`��_���K�%�F�)O�J���-@�R�x�v�����&�A��=����M�:����x�A��� �e�X7׳�-��Eڣ�E�>E��jަlT�/��)@�P��U���	FU}��	"������ZO�l�%�4'�K�`�q�&Xv��z�jP������Y���B��D��M:���2U"R�0~9�#�R��[��ږ������9be��r,cK�3����m�Fq�y;�[[�GbF�4���ۯ8��@�����#_�%y�Jn��DL��yݠ�+
�cKX[F��N�5��*HaP��1�����JrU\�3@���4RZ��W9�%jO:򾕔sˢ�u�uw�Z,��a/b�EU�w+E&���k�yb�Oz@ZlY@��(��LId�[��|%��4ZIXA)ѤRu<8fA�2�O�R
�zҽǫ|�'�Vl�#�G Q�x i�I��"&��x���,Qkm����f��/�'�J��|���VM��]��'�&�p���H>�]�!�ۃ�ԈE���){4�@���D'�~�	�7մDaY��N�j\k5L�~]`�N��n�wG�N��O��f �kns&'�tנ�(�'�@imvĝ�� f��K���q^��Ѧ���VS���AwA�3ُ��$�����ʽ��E�:a;8E.���G�kI�x�ʔ�'ť�}J�����6� ���[���j>�<qZR��P�ӧ�U$�5�� t��P���lg4�3��C�Q��Md�a���8�QM��Q��b����	|zƬ�ۑS#��p�>��DUv�W|?}�e�nb>|�{B+b|�p��؛y^�A�|�u1!�^�8m���ܺ��qº���$�T\W��R�FDϧ�oB%�<�P.a˨�v�M�!�9ة�Ã��َ�r�6�qO;�mC'��O;4o�3:EU�� �B;b����@iY��"'�#�sI[�q'� H���5����3��������N�I'n�U��[V�ٌ ��B����0������\o�?��5SZ���q뫇�F��wA\�BXw��ɪ�.�`��Ϗ���dQ�X��A�ĺv��ݧՇE�v*�ŎE$o����>�`5�~,u�  0&(j/1'޿;
��)^�=?��5�r���,6tҵiֵ9f��A�8o���א|�8���Om��z����RLj![�"�s���ϽC�m������+�Qe���#�զ�ɜha�HK������	�O͜M��翷E���Sk���1��7WL�2&�X�N"��!����hЩ�ƗK��a�vutԐ5�*@b����b"��I��pA��̓��� )�Yi���a"�]�,�m�%��.7U͜a��~$/�B���P<&{!�E:I�D'qr����4��\�����2cdt2�We����[�{����Ъ��p����B+N�c������] Cג�%DPhZd����j���`�_����jsO���Њ�X�:ӻ�x�w�ڲ����������t��uX�}�E������fD�n�"���h�?�?�U?��B�R*�Q����M��vr���?�=�؎�,��dh�)��Ex�.I����nɍjT�{�Agk�^�CD��#1kS�`A�a���H��Ԓ���3���y�M�{!�J��&i�z �M7[�%i��%�=ų�{�脸СJ*��f�c�	��_��s'��eY�0�y!��veC���/��'��A߄�Nf�X�r�:���b�!�Hg��'u�i�c��R�����f��*2��\Q"�2$S�"Q�zФK'xyB�I`�l��uv����u�)�Ո֑!#��y�o,]B����d	�!US�-���\�H��8]>7��t�;mm5���X&T}��4��B0�Y�sl���Y|څ�F�5k�]�%�!���]i� ׎�/fˆ,�y��;�f�>��(������Sȳ��B�J�g�b���.C�ޟ�E���z���]��j��p��֕v�P�7)M�|G$D��X�f���uN��&S~��x�ņ�P����$}�"Z��
�*��OB|k5��)i,�v�����s-U�}�ᔯٮ �yzлxE�;�P���(c&S%�a2�j	��m��J,�2�Ú�[1�:�/�����*k�W�=�#E����(ϧ"OL���S�tԘ;�(�\�{��?u(X)"NlQ6�B+|�7�	`a<bA�D%��b87ݣ�Oa9o�F����t�O��6�z���tdQKY�h�+0���z(IP����C�)ڝ�B]�=�u�)���#��"�]��}�sS�k$3��|8eJ�����AP�K�{�B�yY�7��N�"ۈt4��"�f_�%5��*�R�<��5�!�"F���@�F��G�ϑ��i{��BPhQ��=�����VRBjL�b��E	��%�Wm�a�@j�߬&ip�-g�)Um��1�Lb�_����p�"5����;W�D��4�O)��nn}Ɗ{6Y�#�&�ă���!�@�9�K(��ՙ�: ��M�+,n&��3
�~M��Eخb��C7A}�f���<{)���g'd���KO��>�w:�P��<�'�xw|�8���p77?tsDӬ��Yw�~���#�sq�A/"�g�+�oaOTj��g�;��>xs �ׁ������̬��3�8`?��"����� �!�#B�|	(�b���@ņ��A����H�54ק�gn��6D䵶��$�k�F�ǎ
<���H��]7��;�o�!�W��
��K�N���LY9�����4G�Z�P<�o�SU���µ퐥�� ?�����(- 6a�4U�&���ٷ ���C	2^���Q$h݈�DZ����P���VE}�Jk�u����'rW���o�$���Kb�y5v/'5�hP5[:�u?��$m�"��6��K}B^!	��MX���,ѳ�o u�_R*�9��;�i��#���� Q��m��1���i�.^fl.��Sh�g\�F)��QQ��P��U4��g���"�{����ϩ��D��n1K}m�:���5�cú_�+��S�}P�<��H:�y�����P'p]U7W�is�?��5&��L�S���3Cʇ�"87�?�u�ʐ�?<ƽ�9Y�1���K�2�/u��fb�VH�'t�,R�쭖b
/1�WKz.]p�6+�a�MY��?$(���j��3׃��\��	E��	��d9�)�nvv��C
@��@w����5���qx*H�Y{�#Ef�(+��ƪze�ޫ���5�cxV���ߠ/w/Q,�0������o\i�Y~0:�Ԥ���S�i�쉖,ܑ�-�p�e�F3Հ��)��+�r)���?NQKF�	9P�ք����ó��xaI�D���~`7]�K�D��;�:�w�2���Z��Sy.��Q���}~��vM���/d�xg����v���Y�&��.�`����JD?�����jL����,����"��z�^��jK�Wr�J�"����ϴB��w�����%;��CM�)�-v�e;e*ɰ�j�|5V�=��9���_��0y
�<����.���*�7�?�~x&�34*[w\�� a��r�eJ�������7pu�$��l7�@L�额��6g2���'+��>�"鋭�
��1���y~�%6<"l�3�7�?Fͱ�)½N�F�͙�0���I_����<?��IJ�8O�`�
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(�2���V��Ư3���Z�nm�rķ�I�
��_���������*,4皰c`���(��`l,�uK�����t�!�J~���{�P�*���m���o[��vY�_'�o��#d�4CH�ϳGmɆr8 �~��1m���F�'��,�r�ޮW]�k� ���/�*�tF0"�:
:�}�(�9�E ynf,����b����˥L�:�[�x� N��
�`g��Ya�������;U�\z±�z�"��y��'k<#��ou΅k����k�AY
|����ٽ��7�:D5����؇oUq�~ǘ]gtw�3�����WdX>�_;���Җ&�itn=(���ė��o��C�ߩ���FlA� ��j�����C�����=��'����M)"m������~7��pdu�A|5���?`�9,��Mw8E�Q��˧�~�>����Ɔ��n�LnI���z�C�ݴq�7d�Z�,тT�8�Z˭ ��>����D��әO:ԡ�Љ����!+���	fF4��������-v�bf�G��Ҍ�e��)��'6�֏�?���!Qf�\�ha�i��B��~�P�R�����}�ԫ�Yv��^C�D���f�Mp���Q��ȭ�?gw��1�!y�'I#IO��&�`o� ]�Iq�#���J!�U"0Zǐz�f~�<��a#J�l�}�O����� lk��%�G,�]�[�D��8RYT���������*JA�S�$ �B�(�m��XlxVHYEB    1853     810b�x��:-��W�O5-�C��O܇q��h�-�j�E�_� �:/w*We��.�v��Ta%��W��ʿ�&�1�)�T�V�|پ�}�2��I���"��5�!Y0�U<(��`��v��dh�)��{���Y:�p��c�-����m�B�rp��J���QY�E��YX}���@�v:k���w��q�c����1��>&��X*i����������ש��&�HN�i�k��,�@�7�P}�S?UM��Y� �/�Z�I����?8����ķ��e.����}M�ee�P��z��T��J�k6rF�H��)<���@�ܷ�8��O�MY�Y�|;Zk���m�͏�,�{FE�s��ع*�Y�RNkT,�2�^�^���)|(�N��jM��IC4���oR��˗��&�q��	l��%����&,�����Ѹ
�K}���}P;�P��B֏\�l��;u�R(�� �e7	O�[�Pc��������B���>� ���z��`��9T���՛Q����9��Y��t�Co0��O�(�5��8��ǑHg\���1� -�W� ��<α>��hF�J����#���B~�
x��0�V��q�el��h�L*
���6�KFŪ��E���h��I�eT��@��f��J��v�;[g�ϸ��&���9��4�~-_!�P�Ho��$�2`QʝIi�2��l-]Z�#]
�����p��a當��/P��h�2�X�trv���(��.9�dJ0K�����s�vI��>�c^����]Ex$,��$^�;�\�	�%�`}��)%�7���	�S������D�p�9�f:���麸,��X�#?�2��b���Ǫs������/v��w��h�E&�^�8&eOdkF��EP2��r�Č�D�� ��AG/:�?ZӁY���!�)���{`[��LH�@�(�I�;�	��u��PB��ß�V��l�)������� ~ ���;oP7xpz��=cT_sq�n+_>:7���[��}F�2���z�'�15ph흒��)ܐ�+i���f9#dVJ"�����ݢ���P0I�z��ֻ���{y�ʁ�}ΐ��Oωͽ�13j�5�}=�x�uQù�ix���<�Ev��B&_D��1�A��!l�!�����bz��a���sb&�$/ST+&�Rb"��ݮ�����b@U��c���c�I -��Z0*���A�4�)	©��N�Vv��S/R��<�-+��J�!h`{�$�
�jn�i�ĵ�Kdo����,`���4Z�e��ޮ�>3�߳�_8>�����X��Vi�ԥWpm�b���ݺ�v�!w��p~k���E�Rܰ��{ʦ8
!x�/���^�k������ġ+-s��N
�( J]q�9@Ԋe�}���HĄ,��Z�l�b���oƲIB1A:p!fY���2�\��@���*��!�{�&`*p'�z���(�Z5c.�aI�p [iSp�Ξ�vE�*=�j�0$Ck/�M�|�'.��M�R����ҽ'��s�����PS}Ȏ;Q�M��rh����w��c_����UM��,��V��W[�+%Dl5��fM�^�k� G�����۠��5峕���,G��k;�\~o�R�NI)�絢�rmB�8��ϡ�!��5�%�&���Gy?k�k�n��K�-[�%ա!{�w2�Khp r�w���R�c��_��2|4�F+�4AB�l�8�2
�a{�ViF�IJ��T�q�Lv/�C	�C�ɪ��y�P?�A9�� Z 8��L'<0D��4�7�H�=��פy5���+5�L�Bs�-�?R�_�>��%j�q�t�P�L�́��Ը,=�ի�^�{$�
�Y�@�I�lAn�Xt�6��P�>�4D��T��f`1@U3F�u�����C?v�$[����������ٽJ]9�cmB����ʷ�&�5J
n�ЛZ���Ǟ����:�))[,�Ur$��l�)�t7E}KХ�"c�U��M::�����4
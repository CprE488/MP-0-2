XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R�d��3z�4R�Ú�A����/ho��s?���r��^��s;���)2�%��6�b�b�}i'�����b)PFV�6���ʡ��%ՙ\~4�!�q\教0׊�&��COz�A�<��F�$0���9���<�i,��	���t��'��zW	[/'}����G2q)�@�?��HV�eQ�'zwJj�v��:�u)�`��V�\���,�IE��,
��Ё ,h��Ԥ&��а�kG��Pɟ����]����O�{�eT=��y���V�͋��tAo��]�'�^"��oK(��!c�Y��M|=�bۭI�sE�I�3�x�|�9�}�rVu��(�-�m|�_:]��6����H�N�Jw/H1�Q�+�+�1�<�⦴+�,A�4�N��.��'c����*}�kH�([_�hW���£���9լδQF�E%G�� L���I�^n��zg$$��./.\uA7�܀���Z�H��J��9#͓#����5v��D��J�Y��֠�����{%�Q�+Eivx������ض����&���j��o����;�V%�y�QnsSmU�b���U�J���[�vN����Z2�ng|++7�	�ʶ���(��}���6L;b���tc:u��gJ�*,<�&+�rhqH��{��T�)Wkp'��o����V}��s�T㫦k Q�1�*)<n��l�}�ɳt��	���w}�5B�z� ϑ�b-���WO�+ozY���?��i-XlxVHYEB     f6d     6f0�ڜ�-=��e50����dW���͎?+�0���R��VH*��@ ��+��� m!�rIJ{c�-ZA��m�D�K���dp�'Ϻ��ň�H%�t���{yi�-��t�����q��b0���$^Ӽ[_59��	X¤s��'�m�o��_"N}�c�9����{�B�?�4຀���_�o���)��J�����WbL��-�v�����sM:;���4�O�f���(� ���
h̽��ruJ�*�a�?�e��g���vq�/�M�=/�(��t+e�ef#T��z��[t���;�C�(����`���k6q����5c��7Y���I�Afo:1�D$��*!������%��u��!:V�ӝ[�����dKn�Ĩ��&�r�%Aaɵ��>�<m M|��H�G��~�ډ�?7?ۼ[x����j�(�	:��N�#�Cq�׺'�#�����;�xڢX�&�܂!d�ƫӛ���gJ��X��3����6{��3ƣ�UwT�U��wB�[%��s�w�,x��B� T�4<�Օ�h�[�,n�q�N,���ȚP����m�&�o��v^���?Ճ��,�iEJ:�v�Q������;͞���7����H\*ɼ��'g��e��"�Z�e
1.���Wmt̪�_n��;��>�2�! �{��j���m������Y�W�n�/��O:ke�w<@2�dЄ<�d���UrpF��x`9�\��df!~M�gf����8Т	��}U>əf���s�D ��� �&9�]69@�����0�I��D�|=|��ۉ���r�:�c+�&����[�C�IX�8_%Y҈V�w;�g��]�; ǐ����� ����i��;_�K��7Ax�6�R����M���
����t�>Ť=�L�#-�v7 q��9��P5I��wK��p�q�v�Gu��6�S�Gpm┏�{�����Bj{o�}>y1����xJ��}���9e~ك$��,���!�ƪ�J����l�$h�B����%�P\��/�'\�>P#�X�h������K�Oot�r�tC�	��ڣY*Ii�{ �an���P��/��G�bM���A	��7�S��\Ȑۃ���N���&�X��,	K�6Eߦ.s:|�a�3���^�}T���a׉� &k_���ݍb&y����R'ہ��n�s��K��x�(��*�AB�+~*�!/������l)yRz}.w!�%��j �E�>��b������S$�%��T�-7]
P���Xv�\~�*��K^@���W��F�M�rS����2��c�ӎ4�w��x�;��c�� ����@�pٰ��/[�6mQb��� ��ܪ�zc�~5*��6�8�Ɖ[!P朔����w��?5���"��A_]D�+,kO�1_�J�yT@o�����&OGMi-c�-���8��vDH��`���+��O����SI0Sh��ρ����I}��G׽c�Nf~g��0�D[:3Q�^�.͚���Wp}uI^�L)�Ԍ���G�r�/�ێZ����4�r��ÿ�(wm~N�e����'>�S��|sTLfr�����P�qƎ�(��!�j��HҖX�#��m.{���|*N�6\j����2�c��Kw��P6}�a��A�����
{�p*q��3��*}]�:�h0���<��!�nJ-En,��`��n���"$-��9A�;�ˀ0�����	���)H@ig��6>���7X.]��